module approx_core (
  clk, rst_n, is_random_rsc_dat, is_random_triosy_lz, valid_rsc_dat, valid_triosy_lz,
      epsilon_rsc_dat, epsilon_triosy_lz
);
  input clk;
  input rst_n;
  output is_random_rsc_dat;
  output is_random_triosy_lz;
  output valid_rsc_dat;
  output valid_triosy_lz;
  input epsilon_rsc_dat;
  output epsilon_triosy_lz;


  // Interconnect Declarations
  reg is_random_rsci_idat;
  reg valid_rsci_idat;
  wire epsilon_rsci_idat;
  reg epsilon_triosy_obj_ld;
  wire [4:0] if_4_for_1_acc_tmp;
  wire [5:0] nl_if_4_for_1_acc_tmp;
  wire nand_tmp;
  wire [9:0] if_4_for_mux_50_tmp;
  wire [1:0] mux_3_tmp;
  wire or_2_tmp;
  wire and_dcpl_24;
  wire and_dcpl_25;
  wire and_dcpl_32;
  wire or_dcpl_1;
  wire and_dcpl_39;
  wire and_dcpl_41;
  wire and_dcpl_42;
  wire and_dcpl_43;
  wire or_dcpl_3;
  wire and_dcpl_49;
  wire and_dcpl_59;
  wire and_dcpl_61;
  wire and_dcpl_66;
  wire and_dcpl_67;
  wire or_dcpl_10;
  wire or_dcpl_14;
  wire or_dcpl_20;
  wire or_dcpl_26;
  wire or_dcpl_27;
  wire or_dcpl_28;
  wire or_dcpl_29;
  wire mux_tmp_4;
  wire or_dcpl_33;
  wire or_dcpl_34;
  wire or_dcpl_37;
  wire or_dcpl_43;
  wire or_dcpl_44;
  wire or_dcpl_47;
  wire or_dcpl_54;
  wire or_dcpl_55;
  wire or_dcpl_58;
  wire or_dcpl_65;
  wire or_dcpl_66;
  wire or_dcpl_69;
  wire or_dcpl_76;
  wire or_dcpl_77;
  wire or_dcpl_80;
  wire or_dcpl_81;
  wire or_dcpl_88;
  wire or_dcpl_91;
  wire or_dcpl_98;
  wire or_tmp_12;
  wire or_tmp_14;
  wire mux_tmp_9;
  wire mux_tmp_11;
  wire or_dcpl_100;
  wire or_dcpl_102;
  wire or_dcpl_104;
  wire or_tmp_19;
  wire mux_tmp_16;
  wire or_tmp_21;
  wire and_tmp;
  wire or_tmp_27;
  wire and_tmp_1;
  wire mux_tmp_22;
  wire mux_tmp_23;
  wire mux_tmp_24;
  wire nor_tmp_5;
  wire or_tmp_29;
  wire not_tmp_48;
  wire or_dcpl_118;
  wire or_dcpl_121;
  wire or_dcpl_132;
  wire or_dcpl_139;
  wire or_dcpl_144;
  wire mux_tmp_53;
  wire mux_tmp_57;
  wire or_dcpl_151;
  wire or_dcpl_154;
  wire mux_tmp_61;
  wire or_dcpl_164;
  wire or_dcpl_170;
  wire or_dcpl_174;
  wire or_dcpl_180;
  wire or_dcpl_185;
  wire or_dcpl_188;
  wire if_4_for_and_mdf_sva_1;
  wire exit_if_4_for_lpi_1_dfm_3;
  wire [3:0] j_1_3_0_sva_2;
  wire [4:0] nl_j_1_3_0_sva_2;
  wire exit_if_4_for_lpi_1_dfm_4;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_7_sva_1;
  wire shift_reg_1_sva_0_mx0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_6_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_5_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_4_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_3_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_2_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_1_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_0_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_6_mx0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_5_mx0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_4_mx0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_3_mx0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_2_mx0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_1_mx0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_mx0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_nor_m1c_mx0;
  reg exit_if_4_for_lpi_1_dfm_2;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_1_0_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_1_1_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_1_2_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_1_3_sva_1;
  wire saved_reg_sva_dfm_1_2_mx0;
  wire saved_reg_sva_dfm_1_0_mx0;
  wire saved_reg_sva_dfm_1_1_mx0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_stg_1_3_sva_1;
  reg shift_reg_1_sva_0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_stg_1_2_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_stg_1_1_sva_1;
  reg exitL_exit_if_4_for_2_lpi_1_dfm;
  wire [1:0] skip_sva_dfm_1_0_mx0;
  reg first_sva;
  wire and_91_tmp_1;
  wire [1:0] skip_sva_1_1_0_1;
  wire [2:0] nl_skip_sva_1_1_0_1;
  wire exit_if_4_for_lpi_1_dfm_mx0;
  wire or_psp_mx0;
  wire if_4_for_1_and_stg_1_0_sva_1;
  wire if_4_for_1_and_stg_1_1_sva_1;
  wire if_4_for_1_and_stg_1_2_sva_1;
  wire if_4_for_1_and_stg_1_3_sva_1;
  reg [2:0] j_1_3_0_lpi_1_dfm_2_2_0;
  reg [3:0] j_lpi_1_dfm_1_3_0;
  reg if_4_for_and_mdf_sva_st_1;
  reg mux_1304_itm_1;
  reg [9:0] asn_sft_lpi_1_dfm_st_1;
  reg exitL_exit_approx_sva;
  reg mux_1304_itm_2;
  reg main_stage_0_3;
  reg exitL_exit_if_4_for_2_lpi_1_dfm_st_1_2;
  reg main_stage_0_2;
  reg if_4_for_and_45_itm_1;
  reg operator_24_14_false_AC_TRN_AC_WRAP_1_slc_operator_24_14_false_AC_TRN_AC_WRAP_1_acc_14_svs_1;
  reg shift_reg_1_sva_2;
  reg shift_reg_1_sva_1;
  reg saved_reg_sva_2;
  reg saved_reg_sva_1;
  wire [3:0] j_lpi_1_dfm_3_0_1;
  wire [2:0] j_1_3_0_lpi_1_dfm_2_0_1;
  wire and_55_cse_1;
  wire nor_cse_1;
  reg reg_is_random_triosy_obj_ld_cse;
  wire mux_1368_cse;
  wire mux_1383_cse;
  wire or_247_cse;
  wire nor_47_cse;
  wire or_222_cse;
  wire or_226_cse;
  wire nor_63_cse;
  wire or_99_tmp;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_nor_m1c;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_m1c_3;
  wire or_117_tmp;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_m1c_6;
  wire or_133_tmp;
  wire nor_19_m1c;
  wire or_141_tmp;
  wire nor_20_m1c;
  wire or_152_tmp;
  wire nor_21_m1c;
  wire or_158_tmp;
  wire nor_22_m1c;
  wire or_167_tmp;
  wire nor_23_m1c;
  wire mux_1346_tmp;
  wire nor_24_m1c;
  wire or_183_tmp;
  wire nor_25_m1c;
  wire mux_1353_tmp;
  wire nor_26_m1c;
  wire mux_1313_tmp;
  wire nor_27_m1c;
  wire nand_37_tmp;
  wire nor_28_m1c;
  wire mux_1325_tmp;
  wire nor_29_m1c;
  wire nand_38_tmp;
  wire nor_30_m1c;
  wire or_160_tmp;
  wire nor_31_m1c;
  wire or_170_tmp;
  wire nor_32_m1c;
  wire or_178_tmp;
  wire nor_33_m1c;
  wire or_188_tmp;
  wire nor_34_m1c;
  wire or_251_cse;
  wire mux_1372_cse;
  wire mux_1367_cse;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_nor_3_cse;
  wire if_4_for_and_stg_1_0_sva_1;
  wire if_4_for_and_stg_1_1_sva_1;
  wire if_4_for_and_stg_1_2_sva_1;
  wire if_4_for_and_stg_1_3_sva_1;
  wire [13:0] P1_4_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P1_4_1_23_10_sva_dfm_3;
  wire [13:0] P1_5_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P1_5_1_23_10_sva_dfm_3;
  wire [13:0] P1_1_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P1_1_1_23_10_sva_dfm_3;
  wire [13:0] P1_6_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P1_6_1_23_10_sva_dfm_3;
  wire [13:0] P1_2_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P1_2_1_23_10_sva_dfm_3;
  wire [13:0] P1_7_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P1_7_1_23_10_sva_dfm_3;
  wire [13:0] P1_3_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P1_3_1_23_10_sva_dfm_3;
  wire or_297_tmp;
  wire or_299_tmp;
  wire or_301_tmp;
  wire or_303_tmp;
  wire or_305_tmp;
  wire or_307_tmp;
  wire or_309_tmp;
  wire nand_49_cse;
  wire nand_50_cse;
  wire nand_51_cse;
  wire nand_52_cse;
  wire mux_1310_itm;
  reg [9:0] count_sva;
  wire [10:0] nl_count_sva;
  reg [13:0] P1_3_1_23_10_sva;
  reg [13:0] P1_4_1_23_10_sva;
  reg [13:0] P1_2_1_23_10_sva;
  reg [13:0] P1_5_1_23_10_sva;
  reg [13:0] P1_1_1_23_10_sva;
  reg [13:0] P1_6_1_23_10_sva;
  reg [13:0] P1_7_1_23_10_sva;
  reg [13:0] P2_7_1_23_10_sva;
  reg [13:0] P2_8_1_23_10_sva;
  reg [13:0] P2_6_1_23_10_sva;
  reg [13:0] P2_9_1_23_10_sva;
  reg [13:0] P2_5_1_23_10_sva;
  reg [13:0] P2_10_1_23_10_sva;
  reg [13:0] P2_4_1_23_10_sva;
  reg [13:0] P2_11_1_23_10_sva;
  reg [13:0] P2_3_1_23_10_sva;
  reg [13:0] P2_12_1_23_10_sva;
  reg [13:0] P2_2_1_23_10_sva;
  reg [13:0] P2_13_1_23_10_sva;
  reg [13:0] P2_1_1_23_10_sva;
  reg [13:0] P2_14_1_23_10_sva;
  reg [13:0] P2_0_1_23_10_sva;
  reg [13:0] P2_15_1_23_10_sva;
  reg exit_if_4_for_lpi_1_dfm;
  reg if_4_slc_if_4_acc_1_15_svs;
  reg or_psp;
  reg operator_24_14_false_AC_TRN_AC_WRAP_3_nor_m1c;
  reg operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c;
  reg operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_1;
  reg operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_2;
  reg operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_3;
  reg operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_4;
  reg operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_5;
  reg operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_6;
  reg if_4_for_and_mdf_sva_2;
  reg unequal_tmp_2_1;
  reg unequal_tmp_2_2;
  reg [23:0] sum1_1_lpi_1_dfm_1;
  reg [23:0] sum2_1_lpi_1_dfm_1;
  reg [13:0] operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1;
  reg ln_land_251_lpi_1_dfm_1;
  reg ln_land_252_lpi_1_dfm_1;
  reg ln_if_253_acc_cse_11_sva_1;
  reg ln_and_240_ssc_1;
  reg ln_and_377_ssc_1;
  reg ln_and_242_ssc_1;
  reg ln_and_407_ssc_1;
  reg ln_and_244_ssc_1;
  reg ln_and_379_ssc_1;
  reg ln_and_248_ssc_1;
  reg [13:0] operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1;
  reg ln_1_land_251_lpi_1_dfm_1;
  reg ln_1_land_252_lpi_1_dfm_1;
  reg ln_1_if_253_acc_cse_11_sva_1;
  reg ln_1_and_240_ssc_1;
  reg ln_1_and_377_ssc_1;
  reg ln_1_and_242_ssc_1;
  reg ln_1_and_407_ssc_1;
  reg ln_1_and_244_ssc_1;
  reg ln_1_and_379_ssc_1;
  reg ln_1_and_248_ssc_1;
  reg if_4_slc_if_4_acc_1_15_svs_1;
  reg ln_and_427_itm_1;
  reg ln_1_and_427_itm_1;
  reg [12:0] if_4_aelse_not_itm_1;
  reg saved_reg_sva_0;
  reg ln_ln_mux1h_118_psp_1_12;
  reg ln_ln_mux1h_118_psp_1_11;
  reg ln_ln_mux1h_118_psp_1_10;
  reg ln_ln_mux1h_118_psp_1_8;
  reg ln_ln_mux1h_118_psp_1_7;
  reg ln_ln_mux1h_118_psp_1_6;
  reg ln_ln_mux1h_118_psp_1_5;
  reg ln_ln_mux1h_118_psp_1_4;
  reg ln_ln_mux1h_118_psp_1_3;
  reg ln_ln_mux1h_118_psp_1_2;
  reg ln_ln_mux1h_118_psp_1_1;
  reg ln_ln_mux1h_118_psp_1_0;
  reg ln_1_ln_1_mux1h_118_psp_1_12;
  reg ln_1_ln_1_mux1h_118_psp_1_11;
  reg ln_1_ln_1_mux1h_118_psp_1_10;
  reg ln_1_ln_1_mux1h_118_psp_1_8;
  reg ln_1_ln_1_mux1h_118_psp_1_7;
  reg ln_1_ln_1_mux1h_118_psp_1_6;
  reg ln_1_ln_1_mux1h_118_psp_1_5;
  reg ln_1_ln_1_mux1h_118_psp_1_4;
  reg ln_1_ln_1_mux1h_118_psp_1_3;
  reg ln_1_ln_1_mux1h_118_psp_1_2;
  reg ln_1_ln_1_mux1h_118_psp_1_1;
  reg ln_1_ln_1_mux1h_118_psp_1_0;
  wire ln_land_251_lpi_1_dfm_1_1;
  wire ln_land_252_lpi_1_dfm_1_1;
  wire ln_nor_9_cse_1;
  wire ln_nor_10_cse_1;
  wire ln_and_246_ssc_1;
  wire ln_land_248_lpi_1_dfm_1;
  wire ln_land_249_lpi_1_dfm_1;
  wire ln_land_250_lpi_1_dfm_1;
  wire ln_and_240_ssc_1_1;
  wire ln_land_246_lpi_1_dfm_1;
  wire ln_land_247_lpi_1_dfm_1;
  wire [13:0] operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1;
  wire ln_1_land_251_lpi_1_dfm_1_1;
  wire ln_1_land_252_lpi_1_dfm_1_1;
  wire ln_1_nor_9_cse_1;
  wire ln_1_nor_10_cse_1;
  wire ln_1_and_246_ssc_1;
  wire ln_1_land_248_lpi_1_dfm_1;
  wire ln_1_land_249_lpi_1_dfm_1;
  wire ln_1_land_250_lpi_1_dfm_1;
  wire ln_1_and_240_ssc_1_1;
  wire ln_1_land_246_lpi_1_dfm_1;
  wire ln_1_land_247_lpi_1_dfm_1;
  wire [13:0] operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1;
  wire [14:0] if_4_acc_psp_sva_1;
  wire [15:0] nl_if_4_acc_psp_sva_1;
  wire [23:0] sum1_1_lpi_1_dfm_2_mx0;
  wire [23:0] sum2_1_lpi_1_dfm_1_mx0;
  wire [9:0] asn_sft_lpi_1_dfm_st_1_mx0;
  wire [13:0] P2_0_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P2_8_1_23_10_sva_dfm_1_mx0;
  wire [13:0] operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1;
  wire [14:0] nl_operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1;
  wire [13:0] P2_1_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P2_9_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P2_2_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P2_10_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P2_3_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P2_11_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P2_12_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P2_4_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P2_13_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P2_5_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P2_14_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P2_6_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P2_15_1_23_10_sva_dfm_1_mx0;
  wire [13:0] P2_7_1_23_10_sva_dfm_1_mx0;
  wire [13:0] operator_24_14_false_AC_TRN_AC_WRAP_1_acc_psp_sva_1;
  wire [14:0] nl_operator_24_14_false_AC_TRN_AC_WRAP_1_acc_psp_sva_1;
  wire [13:0] operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1;
  wire [14:0] nl_operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1;
  wire [13:0] operator_24_14_false_AC_TRN_AC_WRAP_3_acc_psp_sva_1;
  wire [14:0] nl_operator_24_14_false_AC_TRN_AC_WRAP_3_acc_psp_sva_1;
  wire [13:0] operator_24_14_false_AC_TRN_AC_WRAP_2_acc_psp_sva_1;
  wire [14:0] nl_operator_24_14_false_AC_TRN_AC_WRAP_2_acc_psp_sva_1;
  wire [13:0] P2_15_2_23_10_sva_mx0;
  wire [13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1;
  wire [14:0] nl_operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1;
  wire [13:0] P2_0_2_23_10_sva_mx0;
  wire [13:0] P2_14_2_23_10_sva_mx0;
  wire [13:0] P2_1_2_23_10_sva_mx0;
  wire [13:0] P2_13_2_23_10_sva_mx0;
  wire [13:0] P2_2_2_23_10_sva_mx0;
  wire [13:0] P2_12_2_23_10_sva_mx0;
  wire [13:0] P2_3_2_23_10_sva_mx0;
  wire [13:0] P2_11_2_23_10_sva_mx0;
  wire [13:0] P2_4_2_23_10_sva_mx0;
  wire [13:0] P2_10_2_23_10_sva_mx0;
  wire [13:0] P2_5_2_23_10_sva_mx0;
  wire [13:0] P2_9_2_23_10_sva_mx0;
  wire [13:0] P2_6_2_23_10_sva_mx0;
  wire [13:0] P2_8_2_23_10_sva_mx0;
  wire [13:0] P2_7_2_23_10_sva_mx0;
  wire [13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1;
  wire [14:0] nl_operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_6_mx0w0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_nor_m1c_mx0w0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_5_mx0w0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_mx0w0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_4_mx0w0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_1_mx0w0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_3_mx0w0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_2_mx0w0;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_11_cse_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_10_cse_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_9_cse_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_8_cse_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_7_cse_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_6_cse_sva_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_4_cse_sva_1;
  wire [13:0] P2_0_1_23_10_sva_dfm_3;
  wire [13:0] P2_1_1_23_10_sva_dfm_3;
  wire [13:0] P2_2_1_23_10_sva_dfm_3;
  wire [13:0] P2_3_1_23_10_sva_dfm_3;
  wire [13:0] P2_4_1_23_10_sva_dfm_3;
  wire [13:0] P2_5_1_23_10_sva_dfm_3;
  wire [13:0] P2_6_1_23_10_sva_dfm_3;
  wire [13:0] P2_7_1_23_10_sva_dfm_3;
  wire [13:0] P2_8_1_23_10_sva_dfm_3;
  wire [13:0] P2_9_1_23_10_sva_dfm_3;
  wire [13:0] P2_10_1_23_10_sva_dfm_3;
  wire [13:0] P2_11_1_23_10_sva_dfm_3;
  wire [13:0] P2_12_1_23_10_sva_dfm_3;
  wire [13:0] P2_13_1_23_10_sva_dfm_3;
  wire [13:0] P2_14_1_23_10_sva_dfm_3;
  wire [13:0] P2_15_1_23_10_sva_dfm_3;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_27_tmp_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_25_tmp_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_23_tmp_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_21_tmp_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_19_tmp_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_17_tmp_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_15_tmp_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_13_tmp_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_12_tmp_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_14_tmp_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_16_tmp_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_18_tmp_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_20_tmp_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_22_tmp_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_24_tmp_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_6_and_26_tmp_1;
  wire and_21_m1c_1;
  wire and_19_m1c_1;
  wire and_17_m1c_1;
  wire and_15_m1c_1;
  wire and_13_m1c_1;
  wire and_11_m1c_1;
  wire and_9_m1c_1;
  wire and_7_m1c_1;
  wire exitL_exit_if_4_for_2_lpi_1_dfm_1;
  wire ln_nor_33_cse_1;
  wire ln_land_17_lpi_1_dfm_1;
  wire ln_land_18_lpi_1_dfm_1;
  wire ln_land_19_lpi_1_dfm_1;
  wire ln_land_20_lpi_1_dfm_1;
  wire ln_land_21_lpi_1_dfm_1;
  wire ln_land_22_lpi_1_dfm_1;
  wire ln_land_23_lpi_1_dfm_1;
  wire ln_land_24_lpi_1_dfm_1;
  wire ln_land_25_lpi_1_dfm_1;
  wire ln_land_26_lpi_1_dfm_1;
  wire ln_land_27_lpi_1_dfm_1;
  wire ln_land_28_lpi_1_dfm_1;
  wire ln_land_29_lpi_1_dfm_1;
  wire ln_land_30_lpi_1_dfm_1;
  wire ln_land_31_lpi_1_dfm_1;
  wire ln_land_32_lpi_1_dfm_1;
  wire ln_land_33_lpi_1_dfm_1;
  wire ln_land_34_lpi_1_dfm_1;
  wire ln_land_35_lpi_1_dfm_1;
  wire ln_land_36_lpi_1_dfm_1;
  wire ln_land_37_lpi_1_dfm_1;
  wire ln_land_38_lpi_1_dfm_1;
  wire ln_land_39_lpi_1_dfm_1;
  wire ln_land_40_lpi_1_dfm_1;
  wire ln_land_41_lpi_1_dfm_1;
  wire ln_land_42_lpi_1_dfm_1;
  wire ln_land_43_lpi_1_dfm_1;
  wire ln_land_44_lpi_1_dfm_1;
  wire ln_land_45_lpi_1_dfm_1;
  wire ln_land_46_lpi_1_dfm_1;
  wire ln_land_47_lpi_1_dfm_1;
  wire ln_land_48_lpi_1_dfm_1;
  wire ln_land_49_lpi_1_dfm_1;
  wire ln_if_50_ln_if_50_and_seb_1;
  wire ln_land_51_lpi_1_dfm_1;
  wire ln_land_52_lpi_1_dfm_1;
  wire ln_land_77_lpi_1_dfm_1;
  wire ln_land_78_lpi_1_dfm_1;
  wire ln_land_79_lpi_1_dfm_1;
  wire ln_land_80_lpi_1_dfm_1;
  wire ln_land_81_lpi_1_dfm_1;
  wire ln_land_82_lpi_1_dfm_1;
  wire ln_land_83_lpi_1_dfm_1;
  wire ln_land_84_lpi_1_dfm_1;
  wire ln_land_85_lpi_1_dfm_1;
  wire ln_land_86_lpi_1_dfm_1;
  wire ln_land_87_lpi_1_dfm_1;
  wire ln_land_88_lpi_1_dfm_1;
  wire ln_land_89_lpi_1_dfm_1;
  wire ln_land_90_lpi_1_dfm_1;
  wire ln_land_91_lpi_1_dfm_1;
  wire ln_land_92_lpi_1_dfm_1;
  wire ln_land_93_lpi_1_dfm_1;
  wire ln_land_94_lpi_1_dfm_1;
  wire ln_land_95_lpi_1_dfm_1;
  wire ln_land_96_lpi_1_dfm_1;
  wire ln_land_97_lpi_1_dfm_1;
  wire ln_land_114_lpi_1_dfm_1;
  wire ln_land_115_lpi_1_dfm_1;
  wire ln_land_116_lpi_1_dfm_1;
  wire ln_land_117_lpi_1_dfm_1;
  wire ln_land_118_lpi_1_dfm_1;
  wire ln_land_119_lpi_1_dfm_1;
  wire ln_land_120_lpi_1_dfm_1;
  wire ln_land_121_lpi_1_dfm_1;
  wire ln_land_122_lpi_1_dfm_1;
  wire ln_land_123_lpi_1_dfm_1;
  wire ln_land_124_lpi_1_dfm_1;
  wire ln_land_125_lpi_1_dfm_1;
  wire ln_land_126_lpi_1_dfm_1;
  wire ln_land_127_lpi_1_dfm_1;
  wire ln_land_128_lpi_1_dfm_1;
  wire ln_land_129_lpi_1_dfm_1;
  wire ln_land_130_lpi_1_dfm_1;
  wire ln_land_131_lpi_1_dfm_1;
  wire ln_land_132_lpi_1_dfm_1;
  wire ln_land_133_lpi_1_dfm_1;
  wire ln_land_134_lpi_1_dfm_1;
  wire ln_land_135_lpi_1_dfm_1;
  wire ln_land_136_lpi_1_dfm_1;
  wire ln_land_137_lpi_1_dfm_1;
  wire ln_land_138_lpi_1_dfm_1;
  wire ln_land_139_lpi_1_dfm_1;
  wire ln_land_140_lpi_1_dfm_1;
  wire ln_and_48_ssc_1;
  wire ln_land_54_lpi_1_dfm_1;
  wire ln_land_55_lpi_1_dfm_1;
  wire ln_land_56_lpi_1_dfm_1;
  wire ln_land_57_lpi_1_dfm_1;
  wire ln_land_58_lpi_1_dfm_1;
  wire ln_land_59_lpi_1_dfm_1;
  wire ln_land_60_lpi_1_dfm_1;
  wire ln_land_61_lpi_1_dfm_1;
  wire ln_land_62_lpi_1_dfm_1;
  wire ln_land_63_lpi_1_dfm_1;
  wire ln_land_64_lpi_1_dfm_1;
  wire ln_land_65_lpi_1_dfm_1;
  wire ln_land_66_lpi_1_dfm_1;
  wire ln_land_67_lpi_1_dfm_1;
  wire ln_land_68_lpi_1_dfm_1;
  wire ln_land_69_lpi_1_dfm_1;
  wire ln_land_70_lpi_1_dfm_1;
  wire ln_land_71_lpi_1_dfm_1;
  wire ln_land_72_lpi_1_dfm_1;
  wire ln_land_73_lpi_1_dfm_1;
  wire ln_land_74_lpi_1_dfm_1;
  wire ln_land_75_lpi_1_dfm_1;
  wire ln_land_76_lpi_1_dfm_1;
  wire ln_land_98_lpi_1_dfm_1;
  wire ln_land_99_lpi_1_dfm_1;
  wire ln_land_100_lpi_1_dfm_1;
  wire ln_land_101_lpi_1_dfm_1;
  wire ln_land_102_lpi_1_dfm_1;
  wire ln_land_103_lpi_1_dfm_1;
  wire ln_land_104_lpi_1_dfm_1;
  wire ln_land_105_lpi_1_dfm_1;
  wire ln_land_106_lpi_1_dfm_1;
  wire ln_land_107_lpi_1_dfm_1;
  wire ln_land_108_lpi_1_dfm_1;
  wire ln_land_109_lpi_1_dfm_1;
  wire ln_land_110_lpi_1_dfm_1;
  wire ln_land_111_lpi_1_dfm_1;
  wire ln_land_112_lpi_1_dfm_1;
  wire ln_land_113_lpi_1_dfm_1;
  wire ln_land_141_lpi_1_dfm_1;
  wire ln_land_142_lpi_1_dfm_1;
  wire ln_and_138_ssc_1;
  wire ln_land_144_lpi_1_dfm_1;
  wire ln_land_172_lpi_1_dfm_1;
  wire ln_land_173_lpi_1_dfm_1;
  wire ln_land_174_lpi_1_dfm_1;
  wire ln_land_175_lpi_1_dfm_1;
  wire ln_land_176_lpi_1_dfm_1;
  wire ln_land_177_lpi_1_dfm_1;
  wire ln_land_178_lpi_1_dfm_1;
  wire ln_land_179_lpi_1_dfm_1;
  wire ln_land_180_lpi_1_dfm_1;
  wire ln_land_181_lpi_1_dfm_1;
  wire ln_land_182_lpi_1_dfm_1;
  wire ln_land_183_lpi_1_dfm_1;
  wire ln_land_184_lpi_1_dfm_1;
  wire ln_land_185_lpi_1_dfm_1;
  wire ln_land_186_lpi_1_dfm_1;
  wire ln_land_187_lpi_1_dfm_1;
  wire ln_land_188_lpi_1_dfm_1;
  wire ln_land_189_lpi_1_dfm_1;
  wire ln_land_190_lpi_1_dfm_1;
  wire ln_land_191_lpi_1_dfm_1;
  wire ln_land_192_lpi_1_dfm_1;
  wire ln_land_193_lpi_1_dfm_1;
  wire ln_land_194_lpi_1_dfm_1;
  wire ln_land_214_lpi_1_dfm_1;
  wire ln_land_215_lpi_1_dfm_1;
  wire ln_land_216_lpi_1_dfm_1;
  wire ln_land_217_lpi_1_dfm_1;
  wire ln_land_218_lpi_1_dfm_1;
  wire ln_land_219_lpi_1_dfm_1;
  wire ln_land_220_lpi_1_dfm_1;
  wire ln_land_221_lpi_1_dfm_1;
  wire ln_land_222_lpi_1_dfm_1;
  wire ln_land_223_lpi_1_dfm_1;
  wire ln_land_224_lpi_1_dfm_1;
  wire ln_land_225_lpi_1_dfm_1;
  wire ln_land_226_lpi_1_dfm_1;
  wire ln_land_227_lpi_1_dfm_1;
  wire ln_land_228_lpi_1_dfm_1;
  wire ln_land_240_lpi_1_dfm_1;
  wire ln_land_241_lpi_1_dfm_1;
  wire ln_land_242_lpi_1_dfm_1;
  wire ln_land_243_lpi_1_dfm_1;
  wire ln_land_244_lpi_1_dfm_1;
  wire ln_and_140_ssc_1;
  wire ln_land_146_lpi_1_dfm_1;
  wire ln_land_147_lpi_1_dfm_1;
  wire ln_land_148_lpi_1_dfm_1;
  wire ln_land_149_lpi_1_dfm_1;
  wire ln_land_150_lpi_1_dfm_1;
  wire ln_land_151_lpi_1_dfm_1;
  wire ln_land_152_lpi_1_dfm_1;
  wire ln_land_153_lpi_1_dfm_1;
  wire ln_land_154_lpi_1_dfm_1;
  wire ln_land_155_lpi_1_dfm_1;
  wire ln_land_156_lpi_1_dfm_1;
  wire ln_land_157_lpi_1_dfm_1;
  wire ln_land_158_lpi_1_dfm_1;
  wire ln_land_159_lpi_1_dfm_1;
  wire ln_land_160_lpi_1_dfm_1;
  wire ln_land_161_lpi_1_dfm_1;
  wire ln_land_162_lpi_1_dfm_1;
  wire ln_land_163_lpi_1_dfm_1;
  wire ln_land_164_lpi_1_dfm_1;
  wire ln_land_165_lpi_1_dfm_1;
  wire ln_land_166_lpi_1_dfm_1;
  wire ln_land_167_lpi_1_dfm_1;
  wire ln_land_168_lpi_1_dfm_1;
  wire ln_land_169_lpi_1_dfm_1;
  wire ln_land_170_lpi_1_dfm_1;
  wire ln_land_171_lpi_1_dfm_1;
  wire ln_land_195_lpi_1_dfm_1;
  wire ln_land_196_lpi_1_dfm_1;
  wire ln_land_197_lpi_1_dfm_1;
  wire ln_land_198_lpi_1_dfm_1;
  wire ln_land_199_lpi_1_dfm_1;
  wire ln_land_200_lpi_1_dfm_1;
  wire ln_land_201_lpi_1_dfm_1;
  wire ln_land_202_lpi_1_dfm_1;
  wire ln_land_203_lpi_1_dfm_1;
  wire ln_land_204_lpi_1_dfm_1;
  wire ln_land_205_lpi_1_dfm_1;
  wire ln_land_206_lpi_1_dfm_1;
  wire ln_land_207_lpi_1_dfm_1;
  wire ln_land_208_lpi_1_dfm_1;
  wire ln_land_209_lpi_1_dfm_1;
  wire ln_land_210_lpi_1_dfm_1;
  wire ln_land_211_lpi_1_dfm_1;
  wire ln_land_212_lpi_1_dfm_1;
  wire ln_land_213_lpi_1_dfm_1;
  wire ln_land_229_lpi_1_dfm_1;
  wire ln_land_230_lpi_1_dfm_1;
  wire ln_land_231_lpi_1_dfm_1;
  wire ln_land_232_lpi_1_dfm_1;
  wire ln_land_233_lpi_1_dfm_1;
  wire ln_land_234_lpi_1_dfm_1;
  wire ln_land_235_lpi_1_dfm_1;
  wire ln_land_236_lpi_1_dfm_1;
  wire ln_land_237_lpi_1_dfm_1;
  wire ln_land_238_lpi_1_dfm_1;
  wire ln_land_239_lpi_1_dfm_1;
  wire ln_nor_3_cse_1;
  wire ln_nor_1_cse_1;
  wire ln_land_8_lpi_1_dfm_1;
  wire ln_land_9_lpi_1_dfm_1;
  wire ln_land_11_lpi_1_dfm_1;
  wire ln_land_13_lpi_1_dfm_1;
  wire ln_land_15_lpi_1_dfm_1;
  wire ln_and_4_ssc_1;
  wire ln_land_10_lpi_1_dfm_1;
  wire ln_land_12_lpi_1_dfm_1;
  wire ln_land_14_lpi_1_dfm_1;
  wire ln_land_16_lpi_1_dfm_1;
  wire ln_and_368_m1c_1;
  wire ln_land_4_lpi_1_dfm_1;
  wire ln_and_2_ssc_1;
  wire ln_land_6_lpi_1_dfm_1;
  wire ln_nor_5_cse_1;
  wire ln_ret_13_0_lpi_1_dfm_258;
  wire ln_land_3_lpi_1_dfm_1;
  wire ln_ln_ln_nor_8_cse_1;
  wire ln_1_nor_33_cse_1;
  wire ln_1_land_17_lpi_1_dfm_1;
  wire ln_1_land_18_lpi_1_dfm_1;
  wire ln_1_land_19_lpi_1_dfm_1;
  wire ln_1_land_20_lpi_1_dfm_1;
  wire ln_1_land_21_lpi_1_dfm_1;
  wire ln_1_land_22_lpi_1_dfm_1;
  wire ln_1_land_23_lpi_1_dfm_1;
  wire ln_1_land_24_lpi_1_dfm_1;
  wire ln_1_land_25_lpi_1_dfm_1;
  wire ln_1_land_26_lpi_1_dfm_1;
  wire ln_1_land_27_lpi_1_dfm_1;
  wire ln_1_land_28_lpi_1_dfm_1;
  wire ln_1_land_29_lpi_1_dfm_1;
  wire ln_1_land_30_lpi_1_dfm_1;
  wire ln_1_land_31_lpi_1_dfm_1;
  wire ln_1_land_32_lpi_1_dfm_1;
  wire ln_1_land_33_lpi_1_dfm_1;
  wire ln_1_land_34_lpi_1_dfm_1;
  wire ln_1_land_35_lpi_1_dfm_1;
  wire ln_1_land_36_lpi_1_dfm_1;
  wire ln_1_land_37_lpi_1_dfm_1;
  wire ln_1_land_38_lpi_1_dfm_1;
  wire ln_1_land_39_lpi_1_dfm_1;
  wire ln_1_land_40_lpi_1_dfm_1;
  wire ln_1_land_41_lpi_1_dfm_1;
  wire ln_1_land_42_lpi_1_dfm_1;
  wire ln_1_land_43_lpi_1_dfm_1;
  wire ln_1_land_44_lpi_1_dfm_1;
  wire ln_1_land_45_lpi_1_dfm_1;
  wire ln_1_land_46_lpi_1_dfm_1;
  wire ln_1_land_47_lpi_1_dfm_1;
  wire ln_1_land_48_lpi_1_dfm_1;
  wire ln_1_land_49_lpi_1_dfm_1;
  wire ln_1_if_50_ln_1_if_50_and_seb_1;
  wire ln_1_land_51_lpi_1_dfm_1;
  wire ln_1_land_52_lpi_1_dfm_1;
  wire ln_1_land_77_lpi_1_dfm_1;
  wire ln_1_land_78_lpi_1_dfm_1;
  wire ln_1_land_79_lpi_1_dfm_1;
  wire ln_1_land_80_lpi_1_dfm_1;
  wire ln_1_land_81_lpi_1_dfm_1;
  wire ln_1_land_82_lpi_1_dfm_1;
  wire ln_1_land_83_lpi_1_dfm_1;
  wire ln_1_land_84_lpi_1_dfm_1;
  wire ln_1_land_85_lpi_1_dfm_1;
  wire ln_1_land_86_lpi_1_dfm_1;
  wire ln_1_land_87_lpi_1_dfm_1;
  wire ln_1_land_88_lpi_1_dfm_1;
  wire ln_1_land_89_lpi_1_dfm_1;
  wire ln_1_land_90_lpi_1_dfm_1;
  wire ln_1_land_91_lpi_1_dfm_1;
  wire ln_1_land_92_lpi_1_dfm_1;
  wire ln_1_land_93_lpi_1_dfm_1;
  wire ln_1_land_94_lpi_1_dfm_1;
  wire ln_1_land_95_lpi_1_dfm_1;
  wire ln_1_land_96_lpi_1_dfm_1;
  wire ln_1_land_97_lpi_1_dfm_1;
  wire ln_1_land_114_lpi_1_dfm_1;
  wire ln_1_land_115_lpi_1_dfm_1;
  wire ln_1_land_116_lpi_1_dfm_1;
  wire ln_1_land_117_lpi_1_dfm_1;
  wire ln_1_land_118_lpi_1_dfm_1;
  wire ln_1_land_119_lpi_1_dfm_1;
  wire ln_1_land_120_lpi_1_dfm_1;
  wire ln_1_land_121_lpi_1_dfm_1;
  wire ln_1_land_122_lpi_1_dfm_1;
  wire ln_1_land_123_lpi_1_dfm_1;
  wire ln_1_land_124_lpi_1_dfm_1;
  wire ln_1_land_125_lpi_1_dfm_1;
  wire ln_1_land_126_lpi_1_dfm_1;
  wire ln_1_land_127_lpi_1_dfm_1;
  wire ln_1_land_128_lpi_1_dfm_1;
  wire ln_1_land_129_lpi_1_dfm_1;
  wire ln_1_land_130_lpi_1_dfm_1;
  wire ln_1_land_131_lpi_1_dfm_1;
  wire ln_1_land_132_lpi_1_dfm_1;
  wire ln_1_land_133_lpi_1_dfm_1;
  wire ln_1_land_134_lpi_1_dfm_1;
  wire ln_1_land_135_lpi_1_dfm_1;
  wire ln_1_land_136_lpi_1_dfm_1;
  wire ln_1_land_137_lpi_1_dfm_1;
  wire ln_1_land_138_lpi_1_dfm_1;
  wire ln_1_land_139_lpi_1_dfm_1;
  wire ln_1_land_140_lpi_1_dfm_1;
  wire ln_1_and_48_ssc_1;
  wire ln_1_land_54_lpi_1_dfm_1;
  wire ln_1_land_55_lpi_1_dfm_1;
  wire ln_1_land_56_lpi_1_dfm_1;
  wire ln_1_land_57_lpi_1_dfm_1;
  wire ln_1_land_58_lpi_1_dfm_1;
  wire ln_1_land_59_lpi_1_dfm_1;
  wire ln_1_land_60_lpi_1_dfm_1;
  wire ln_1_land_61_lpi_1_dfm_1;
  wire ln_1_land_62_lpi_1_dfm_1;
  wire ln_1_land_63_lpi_1_dfm_1;
  wire ln_1_land_64_lpi_1_dfm_1;
  wire ln_1_land_65_lpi_1_dfm_1;
  wire ln_1_land_66_lpi_1_dfm_1;
  wire ln_1_land_67_lpi_1_dfm_1;
  wire ln_1_land_68_lpi_1_dfm_1;
  wire ln_1_land_69_lpi_1_dfm_1;
  wire ln_1_land_70_lpi_1_dfm_1;
  wire ln_1_land_71_lpi_1_dfm_1;
  wire ln_1_land_72_lpi_1_dfm_1;
  wire ln_1_land_73_lpi_1_dfm_1;
  wire ln_1_land_74_lpi_1_dfm_1;
  wire ln_1_land_75_lpi_1_dfm_1;
  wire ln_1_land_76_lpi_1_dfm_1;
  wire ln_1_land_98_lpi_1_dfm_1;
  wire ln_1_land_99_lpi_1_dfm_1;
  wire ln_1_land_100_lpi_1_dfm_1;
  wire ln_1_land_101_lpi_1_dfm_1;
  wire ln_1_land_102_lpi_1_dfm_1;
  wire ln_1_land_103_lpi_1_dfm_1;
  wire ln_1_land_104_lpi_1_dfm_1;
  wire ln_1_land_105_lpi_1_dfm_1;
  wire ln_1_land_106_lpi_1_dfm_1;
  wire ln_1_land_107_lpi_1_dfm_1;
  wire ln_1_land_108_lpi_1_dfm_1;
  wire ln_1_land_109_lpi_1_dfm_1;
  wire ln_1_land_110_lpi_1_dfm_1;
  wire ln_1_land_111_lpi_1_dfm_1;
  wire ln_1_land_112_lpi_1_dfm_1;
  wire ln_1_land_113_lpi_1_dfm_1;
  wire ln_1_land_141_lpi_1_dfm_1;
  wire ln_1_land_142_lpi_1_dfm_1;
  wire ln_1_and_138_ssc_1;
  wire ln_1_land_144_lpi_1_dfm_1;
  wire ln_1_land_172_lpi_1_dfm_1;
  wire ln_1_land_173_lpi_1_dfm_1;
  wire ln_1_land_174_lpi_1_dfm_1;
  wire ln_1_land_175_lpi_1_dfm_1;
  wire ln_1_land_176_lpi_1_dfm_1;
  wire ln_1_land_177_lpi_1_dfm_1;
  wire ln_1_land_178_lpi_1_dfm_1;
  wire ln_1_land_179_lpi_1_dfm_1;
  wire ln_1_land_180_lpi_1_dfm_1;
  wire ln_1_land_181_lpi_1_dfm_1;
  wire ln_1_land_182_lpi_1_dfm_1;
  wire ln_1_land_183_lpi_1_dfm_1;
  wire ln_1_land_184_lpi_1_dfm_1;
  wire ln_1_land_185_lpi_1_dfm_1;
  wire ln_1_land_186_lpi_1_dfm_1;
  wire ln_1_land_187_lpi_1_dfm_1;
  wire ln_1_land_188_lpi_1_dfm_1;
  wire ln_1_land_189_lpi_1_dfm_1;
  wire ln_1_land_190_lpi_1_dfm_1;
  wire ln_1_land_191_lpi_1_dfm_1;
  wire ln_1_land_192_lpi_1_dfm_1;
  wire ln_1_land_193_lpi_1_dfm_1;
  wire ln_1_land_194_lpi_1_dfm_1;
  wire ln_1_land_214_lpi_1_dfm_1;
  wire ln_1_land_215_lpi_1_dfm_1;
  wire ln_1_land_216_lpi_1_dfm_1;
  wire ln_1_land_217_lpi_1_dfm_1;
  wire ln_1_land_218_lpi_1_dfm_1;
  wire ln_1_land_219_lpi_1_dfm_1;
  wire ln_1_land_220_lpi_1_dfm_1;
  wire ln_1_land_221_lpi_1_dfm_1;
  wire ln_1_land_222_lpi_1_dfm_1;
  wire ln_1_land_223_lpi_1_dfm_1;
  wire ln_1_land_224_lpi_1_dfm_1;
  wire ln_1_land_225_lpi_1_dfm_1;
  wire ln_1_land_226_lpi_1_dfm_1;
  wire ln_1_land_227_lpi_1_dfm_1;
  wire ln_1_land_228_lpi_1_dfm_1;
  wire ln_1_land_240_lpi_1_dfm_1;
  wire ln_1_land_241_lpi_1_dfm_1;
  wire ln_1_land_242_lpi_1_dfm_1;
  wire ln_1_land_243_lpi_1_dfm_1;
  wire ln_1_land_244_lpi_1_dfm_1;
  wire ln_1_and_140_ssc_1;
  wire ln_1_land_146_lpi_1_dfm_1;
  wire ln_1_land_147_lpi_1_dfm_1;
  wire ln_1_land_148_lpi_1_dfm_1;
  wire ln_1_land_149_lpi_1_dfm_1;
  wire ln_1_land_150_lpi_1_dfm_1;
  wire ln_1_land_151_lpi_1_dfm_1;
  wire ln_1_land_152_lpi_1_dfm_1;
  wire ln_1_land_153_lpi_1_dfm_1;
  wire ln_1_land_154_lpi_1_dfm_1;
  wire ln_1_land_155_lpi_1_dfm_1;
  wire ln_1_land_156_lpi_1_dfm_1;
  wire ln_1_land_157_lpi_1_dfm_1;
  wire ln_1_land_158_lpi_1_dfm_1;
  wire ln_1_land_159_lpi_1_dfm_1;
  wire ln_1_land_160_lpi_1_dfm_1;
  wire ln_1_land_161_lpi_1_dfm_1;
  wire ln_1_land_162_lpi_1_dfm_1;
  wire ln_1_land_163_lpi_1_dfm_1;
  wire ln_1_land_164_lpi_1_dfm_1;
  wire ln_1_land_165_lpi_1_dfm_1;
  wire ln_1_land_166_lpi_1_dfm_1;
  wire ln_1_land_167_lpi_1_dfm_1;
  wire ln_1_land_168_lpi_1_dfm_1;
  wire ln_1_land_169_lpi_1_dfm_1;
  wire ln_1_land_170_lpi_1_dfm_1;
  wire ln_1_land_171_lpi_1_dfm_1;
  wire ln_1_land_195_lpi_1_dfm_1;
  wire ln_1_land_196_lpi_1_dfm_1;
  wire ln_1_land_197_lpi_1_dfm_1;
  wire ln_1_land_198_lpi_1_dfm_1;
  wire ln_1_land_199_lpi_1_dfm_1;
  wire ln_1_land_200_lpi_1_dfm_1;
  wire ln_1_land_201_lpi_1_dfm_1;
  wire ln_1_land_202_lpi_1_dfm_1;
  wire ln_1_land_203_lpi_1_dfm_1;
  wire ln_1_land_204_lpi_1_dfm_1;
  wire ln_1_land_205_lpi_1_dfm_1;
  wire ln_1_land_206_lpi_1_dfm_1;
  wire ln_1_land_207_lpi_1_dfm_1;
  wire ln_1_land_208_lpi_1_dfm_1;
  wire ln_1_land_209_lpi_1_dfm_1;
  wire ln_1_land_210_lpi_1_dfm_1;
  wire ln_1_land_211_lpi_1_dfm_1;
  wire ln_1_land_212_lpi_1_dfm_1;
  wire ln_1_land_213_lpi_1_dfm_1;
  wire ln_1_land_229_lpi_1_dfm_1;
  wire ln_1_land_230_lpi_1_dfm_1;
  wire ln_1_land_231_lpi_1_dfm_1;
  wire ln_1_land_232_lpi_1_dfm_1;
  wire ln_1_land_233_lpi_1_dfm_1;
  wire ln_1_land_234_lpi_1_dfm_1;
  wire ln_1_land_235_lpi_1_dfm_1;
  wire ln_1_land_236_lpi_1_dfm_1;
  wire ln_1_land_237_lpi_1_dfm_1;
  wire ln_1_land_238_lpi_1_dfm_1;
  wire ln_1_land_239_lpi_1_dfm_1;
  wire ln_1_nor_3_cse_1;
  wire ln_1_nor_1_cse_1;
  wire ln_1_land_8_lpi_1_dfm_1;
  wire ln_1_land_9_lpi_1_dfm_1;
  wire ln_1_land_11_lpi_1_dfm_1;
  wire ln_1_land_13_lpi_1_dfm_1;
  wire ln_1_land_15_lpi_1_dfm_1;
  wire ln_1_and_4_ssc_1;
  wire ln_1_land_10_lpi_1_dfm_1;
  wire ln_1_land_12_lpi_1_dfm_1;
  wire ln_1_land_14_lpi_1_dfm_1;
  wire ln_1_land_16_lpi_1_dfm_1;
  wire ln_1_and_368_m1c_1;
  wire ln_1_land_4_lpi_1_dfm_1;
  wire ln_1_and_2_ssc_1;
  wire ln_1_land_6_lpi_1_dfm_1;
  wire ln_1_nor_5_cse_1;
  wire ln_1_ret_13_0_lpi_1_dfm_257;
  wire ln_1_land_3_lpi_1_dfm_1;
  wire ln_1_ln_1_ln_1_nor_8_cse_1;
  wire if_4_for_1_and_stg_2_7_sva_1;
  wire if_4_for_1_and_stg_2_0_sva_1;
  wire if_4_for_1_and_stg_2_6_sva_1;
  wire if_4_for_1_and_stg_2_1_sva_1;
  wire if_4_for_1_and_stg_2_5_sva_1;
  wire if_4_for_1_and_stg_2_2_sva_1;
  wire if_4_for_1_and_stg_2_4_sva_1;
  wire if_4_for_1_and_stg_2_3_sva_1;
  wire skip_static_init_or_ssc;
  reg reg_skip_ftd;
  reg [1:0] reg_skip_ftd_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_38_cse;
  wire or_tmp_82;
  wire or_tmp_83;
  wire or_tmp_85;
  wire not_tmp_87;
  wire or_tmp_86;
  wire mux_tmp_96;
  wire or_tmp_88;
  wire or_tmp_89;
  wire or_tmp_90;
  wire not_tmp_88;
  wire mux_tmp_104;
  wire mux_tmp_105;
  wire or_tmp_93;
  wire mux_tmp_113;
  wire not_tmp_91;
  wire or_tmp_100;
  wire not_tmp_92;
  wire or_tmp_101;
  wire mux_tmp_119;
  wire or_tmp_104;
  wire mux_tmp_122;
  wire or_tmp_105;
  wire mux_tmp_125;
  wire mux_tmp_126;
  wire mux_tmp_130;
  wire mux_tmp_136;
  wire mux_tmp_141;
  wire mux_tmp_143;
  wire mux_tmp_145;
  wire or_tmp_121;
  wire or_tmp_125;
  wire not_tmp_104;
  wire or_tmp_127;
  wire mux_tmp_156;
  wire or_tmp_129;
  wire or_tmp_131;
  wire mux_tmp_157;
  wire or_tmp_133;
  wire nand_tmp_13;
  wire mux_tmp_162;
  wire mux_tmp_167;
  wire or_tmp_143;
  wire mux_tmp_172;
  wire or_tmp_146;
  wire mux_tmp_173;
  wire mux_tmp_174;
  wire mux_tmp_177;
  wire mux_tmp_183;
  wire mux_tmp_186;
  wire mux_tmp_193;
  wire nor_tmp_32;
  wire mux_tmp_198;
  wire not_tmp_120;
  wire mux_tmp_199;
  wire or_tmp_161;
  wire mux_tmp_200;
  wire nor_tmp_35;
  wire mux_tmp_205;
  wire mux_tmp_208;
  wire mux_tmp_211;
  wire mux_tmp_213;
  wire not_tmp_127;
  wire not_tmp_131;
  wire or_tmp_170;
  wire not_tmp_135;
  wire mux_tmp_228;
  wire or_tmp_176;
  wire mux_tmp_233;
  wire mux_tmp_235;
  wire mux_tmp_237;
  wire mux_tmp_240;
  wire nand_tmp_16;
  wire mux_tmp_251;
  wire or_tmp_186;
  wire or_tmp_187;
  wire mux_tmp_256;
  wire or_tmp_190;
  wire mux_tmp_259;
  wire mux_tmp_264;
  wire mux_tmp_265;
  wire mux_tmp_268;
  wire mux_tmp_279;
  wire or_tmp_205;
  wire mux_tmp_284;
  wire mux_tmp_285;
  wire or_tmp_209;
  wire or_tmp_210;
  wire mux_tmp_286;
  wire mux_tmp_291;
  wire mux_tmp_294;
  wire or_tmp_216;
  wire not_tmp_151;
  wire mux_tmp_298;
  wire mux_tmp_308;
  wire or_tmp_227;
  wire not_tmp_154;
  wire mux_tmp_314;
  wire or_tmp_229;
  wire or_tmp_231;
  wire mux_tmp_317;
  wire mux_tmp_319;
  wire nor_tmp_52;
  wire not_tmp_160;
  wire mux_tmp_326;
  wire mux_tmp_330;
  wire and_tmp_12;
  wire mux_tmp_339;
  wire or_tmp_240;
  wire mux_tmp_346;
  wire or_tmp_245;
  wire or_tmp_248;
  wire and_tmp_13;
  wire mux_tmp_350;
  wire mux_tmp_356;
  wire mux_tmp_361;
  wire mux_tmp_362;
  wire nand_tmp_19;
  wire not_tmp_175;
  wire mux_tmp_366;
  wire mux_tmp_378;
  wire or_tmp_269;
  wire nand_tmp_20;
  wire mux_tmp_385;
  wire mux_tmp_387;
  wire mux_tmp_390;
  wire mux_tmp_394;
  wire mux_tmp_395;
  wire mux_tmp_401;
  wire not_tmp_188;
  wire mux_tmp_408;
  wire mux_tmp_410;
  wire or_tmp_294;
  wire nor_tmp_78;
  wire mux_tmp_416;
  wire nor_tmp_80;
  wire mux_tmp_422;
  wire not_tmp_199;
  wire mux_tmp_425;
  wire mux_tmp_433;
  wire mux_tmp_440;
  wire or_tmp_306;
  wire mux_tmp_444;
  wire or_tmp_308;
  wire or_tmp_309;
  wire or_tmp_310;
  wire and_tmp_15;
  wire or_tmp_323;
  wire or_tmp_325;
  wire mux_tmp_467;
  wire or_tmp_329;
  wire or_tmp_334;
  wire mux_tmp_479;
  wire mux_tmp_480;
  wire or_tmp_336;
  wire mux_tmp_485;
  wire mux_tmp_486;
  wire mux_tmp_487;
  wire mux_tmp_497;
  wire mux_tmp_498;
  wire or_tmp_343;
  wire or_tmp_346;
  wire mux_tmp_503;
  wire or_tmp_347;
  wire mux_tmp_509;
  wire and_tmp_17;
  wire mux_tmp_524;
  wire or_tmp_356;
  wire or_tmp_357;
  wire nor_tmp_112;
  wire mux_tmp_533;
  wire mux_tmp_534;
  wire mux_tmp_538;
  wire not_tmp_236;
  wire mux_tmp_546;
  wire nor_tmp_119;
  wire mux_tmp_549;
  wire nand_tmp_28;
  wire or_tmp_370;
  wire and_276_cse;
  wire or_325_cse;
  wire or_324_cse;
  wire nand_101_cse;
  wire nor_149_cse;
  wire nor_159_cse;
  wire nand_112_cse;
  wire and_294_cse;
  wire nand_128_cse;
  wire nand_116_cse;
  wire or_482_cse;
  wire nand_125_cse;
  wire and_317_cse;
  wire and_351_cse;
  wire and_298_cse;
  wire nor_87_cse;
  wire or_446_cse;
  wire mux_1558_cse;
  wire or_341_cse;
  wire or_387_cse;
  wire or_327_cse;
  wire mux_1756_cse;
  wire nand_150_cse;
  wire or_546_cse;
  wire mux_1547_cse;
  wire nand_86_cse;
  wire if_4_acc_1_itm_15_1;
  wire ln_if_253_acc_itm_11_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_acc_itm_14_1;
  wire ln_1_if_253_acc_itm_11_1;
  wire operator_24_14_false_AC_TRN_AC_WRAP_1_acc_itm_14_1;
  wire ln_if_252_acc_itm_12_1;
  wire ln_if_244_acc_itm_14_1;
  wire ln_if_245_acc_itm_13_1;
  wire ln_if_251_acc_itm_10_1;
  wire ln_if_250_acc_itm_12_1;
  wire ln_if_249_acc_itm_11_1;
  wire ln_if_248_acc_itm_12_1;
  wire ln_if_247_acc_itm_9_1;
  wire ln_if_246_acc_itm_14_1;
  wire ln_if_144_acc_itm_14_1;
  wire ln_if_145_acc_itm_13_1;
  wire ln_if_243_acc_itm_12_1;
  wire ln_if_242_acc_itm_14_1;
  wire ln_if_241_acc_itm_13_1;
  wire ln_if_240_acc_itm_14_1;
  wire ln_if_239_acc_itm_11_1;
  wire ln_if_238_acc_itm_14_1;
  wire ln_if_237_acc_itm_13_1;
  wire ln_if_236_acc_itm_14_1;
  wire ln_if_235_acc_itm_12_1;
  wire ln_if_234_acc_itm_14_1;
  wire ln_if_233_acc_itm_13_1;
  wire ln_if_232_acc_itm_14_1;
  wire ln_if_231_acc_itm_10_1;
  wire ln_if_230_acc_itm_14_1;
  wire ln_if_229_acc_itm_13_1;
  wire ln_if_228_acc_itm_14_1;
  wire ln_if_227_acc_itm_12_1;
  wire ln_if_226_acc_itm_14_1;
  wire ln_if_225_acc_itm_13_1;
  wire ln_if_224_acc_itm_14_1;
  wire ln_if_223_acc_itm_11_1;
  wire ln_if_222_acc_itm_14_1;
  wire ln_if_221_acc_itm_13_1;
  wire ln_if_220_acc_itm_14_1;
  wire ln_if_219_acc_itm_12_1;
  wire ln_if_218_acc_itm_14_1;
  wire ln_if_217_acc_itm_13_1;
  wire ln_if_216_acc_itm_14_1;
  wire ln_if_215_acc_itm_8_1;
  wire ln_if_214_acc_itm_14_1;
  wire ln_if_213_acc_itm_13_1;
  wire ln_if_212_acc_itm_14_1;
  wire ln_if_211_acc_itm_12_1;
  wire ln_if_210_acc_itm_14_1;
  wire ln_if_209_acc_itm_13_1;
  wire ln_if_208_acc_itm_14_1;
  wire ln_if_207_acc_itm_11_1;
  wire ln_if_206_acc_itm_14_1;
  wire ln_if_205_acc_itm_13_1;
  wire ln_if_204_acc_itm_14_1;
  wire ln_if_203_acc_itm_12_1;
  wire ln_if_202_acc_itm_14_1;
  wire ln_if_201_acc_itm_13_1;
  wire ln_if_200_acc_itm_14_1;
  wire ln_if_199_acc_itm_10_1;
  wire ln_if_198_acc_itm_14_1;
  wire ln_if_197_acc_itm_13_1;
  wire ln_if_196_acc_itm_14_1;
  wire ln_if_195_acc_itm_12_1;
  wire ln_if_194_acc_itm_14_1;
  wire ln_if_193_acc_itm_13_1;
  wire ln_if_192_acc_itm_14_1;
  wire ln_if_191_acc_itm_11_1;
  wire ln_if_190_acc_itm_14_1;
  wire ln_if_189_acc_itm_13_1;
  wire ln_if_188_acc_itm_14_1;
  wire ln_if_187_acc_itm_12_1;
  wire ln_if_186_acc_itm_14_1;
  wire ln_if_185_acc_itm_13_1;
  wire ln_if_184_acc_itm_14_1;
  wire ln_if_183_acc_itm_9_1;
  wire ln_if_182_acc_itm_14_1;
  wire ln_if_181_acc_itm_13_1;
  wire ln_if_180_acc_itm_14_1;
  wire ln_if_179_acc_itm_12_1;
  wire ln_if_178_acc_itm_14_1;
  wire ln_if_177_acc_itm_13_1;
  wire ln_if_176_acc_itm_14_1;
  wire ln_if_175_acc_itm_11_1;
  wire ln_if_174_acc_itm_14_1;
  wire ln_if_173_acc_itm_13_1;
  wire ln_if_172_acc_itm_14_1;
  wire ln_if_171_acc_itm_12_1;
  wire ln_if_170_acc_itm_14_1;
  wire ln_if_169_acc_itm_13_1;
  wire ln_if_168_acc_itm_14_1;
  wire ln_if_167_acc_itm_10_1;
  wire ln_if_166_acc_itm_14_1;
  wire ln_if_165_acc_itm_13_1;
  wire ln_if_164_acc_itm_14_1;
  wire ln_if_163_acc_itm_12_1;
  wire ln_if_162_acc_itm_14_1;
  wire ln_if_161_acc_itm_13_1;
  wire ln_if_160_acc_itm_14_1;
  wire ln_if_159_acc_itm_11_1;
  wire ln_if_158_acc_itm_14_1;
  wire ln_if_157_acc_itm_13_1;
  wire ln_if_156_acc_itm_14_1;
  wire ln_if_155_acc_itm_12_1;
  wire ln_if_154_acc_itm_14_1;
  wire ln_if_153_acc_itm_13_1;
  wire ln_if_152_acc_itm_14_1;
  wire ln_if_151_acc_itm_7_1;
  wire ln_if_150_acc_itm_14_1;
  wire ln_if_149_acc_itm_13_1;
  wire ln_if_148_acc_itm_14_1;
  wire ln_if_147_acc_itm_12_1;
  wire ln_if_146_acc_itm_14_1;
  wire ln_if_142_acc_itm_14_1;
  wire ln_if_143_acc_itm_11_1;
  wire ln_if_141_acc_itm_13_1;
  wire ln_if_140_acc_itm_14_1;
  wire ln_if_52_acc_itm_14_1;
  wire ln_if_53_acc_itm_14_1;
  wire ln_if_49_acc_itm_12_1;
  wire ln_if_50_acc_itm_14_1;
  wire ln_if_6_acc_itm_8_1;
  wire ln_if_7_acc_itm_5_1;
  wire ln_if_139_acc_itm_12_1;
  wire ln_if_138_acc_itm_14_1;
  wire ln_if_137_acc_itm_13_1;
  wire ln_if_136_acc_itm_14_1;
  wire ln_if_135_acc_itm_10_1;
  wire ln_if_134_acc_itm_14_1;
  wire ln_if_133_acc_itm_13_1;
  wire ln_if_132_acc_itm_14_1;
  wire ln_if_131_acc_itm_12_1;
  wire ln_if_130_acc_itm_14_1;
  wire ln_if_129_acc_itm_13_1;
  wire ln_if_128_acc_itm_14_1;
  wire ln_if_127_acc_itm_11_1;
  wire ln_if_126_acc_itm_14_1;
  wire ln_if_125_acc_itm_13_1;
  wire ln_if_124_acc_itm_14_1;
  wire ln_if_123_acc_itm_12_1;
  wire ln_if_122_acc_itm_14_1;
  wire ln_if_121_acc_itm_13_1;
  wire ln_if_120_acc_itm_14_1;
  wire ln_if_119_acc_itm_9_1;
  wire ln_if_118_acc_itm_14_1;
  wire ln_if_117_acc_itm_13_1;
  wire ln_if_116_acc_itm_14_1;
  wire ln_if_115_acc_itm_14_1;
  wire ln_if_114_acc_itm_10_1;
  wire ln_if_113_acc_itm_14_1;
  wire ln_if_112_acc_itm_13_1;
  wire ln_if_111_acc_itm_14_1;
  wire ln_if_110_acc_itm_12_1;
  wire ln_if_109_acc_itm_14_1;
  wire ln_if_108_acc_itm_14_1;
  wire ln_if_107_acc_itm_13_1;
  wire ln_if_106_acc_itm_14_1;
  wire ln_if_105_acc_itm_12_1;
  wire ln_if_104_acc_itm_14_1;
  wire ln_if_103_acc_itm_13_1;
  wire ln_if_102_acc_itm_14_1;
  wire ln_if_101_acc_itm_14_1;
  wire ln_if_100_acc_itm_12_1;
  wire ln_if_99_acc_itm_14_1;
  wire ln_if_98_acc_itm_13_1;
  wire ln_if_97_acc_itm_14_1;
  wire ln_if_96_acc_itm_11_1;
  wire ln_if_95_acc_itm_14_1;
  wire ln_if_94_acc_itm_14_1;
  wire ln_if_93_acc_itm_13_1;
  wire ln_if_92_acc_itm_14_1;
  wire ln_if_91_acc_itm_11_1;
  wire ln_if_90_acc_itm_14_1;
  wire ln_if_89_acc_itm_13_1;
  wire ln_if_88_acc_itm_14_1;
  wire ln_if_87_acc_itm_14_1;
  wire ln_if_86_acc_itm_11_1;
  wire ln_if_85_acc_itm_14_1;
  wire ln_if_84_acc_itm_13_1;
  wire ln_if_83_acc_itm_14_1;
  wire ln_if_82_acc_itm_12_1;
  wire ln_if_81_acc_itm_14_1;
  wire ln_if_80_acc_itm_14_1;
  wire ln_if_79_acc_itm_13_1;
  wire ln_if_78_acc_itm_14_1;
  wire ln_if_77_acc_itm_12_1;
  wire ln_if_76_acc_itm_14_1;
  wire ln_if_75_acc_itm_13_1;
  wire ln_if_74_acc_itm_14_1;
  wire ln_if_73_acc_itm_14_1;
  wire ln_if_72_acc_itm_12_1;
  wire ln_if_71_acc_itm_14_1;
  wire ln_if_70_acc_itm_13_1;
  wire ln_if_69_acc_itm_14_1;
  wire ln_if_68_acc_itm_8_1;
  wire ln_if_67_acc_itm_14_1;
  wire ln_if_66_acc_itm_14_1;
  wire ln_if_65_acc_itm_13_1;
  wire ln_if_64_acc_itm_14_1;
  wire ln_if_63_acc_itm_10_1;
  wire ln_if_62_acc_itm_14_1;
  wire ln_if_61_acc_itm_13_1;
  wire ln_if_60_acc_itm_14_1;
  wire ln_if_59_acc_itm_14_1;
  wire ln_if_58_acc_itm_9_1;
  wire ln_if_57_acc_itm_14_1;
  wire ln_if_56_acc_itm_13_1;
  wire ln_if_55_acc_itm_14_1;
  wire ln_if_54_acc_itm_12_1;
  wire ln_if_51_acc_itm_13_1;
  wire ln_if_48_acc_itm_14_1;
  wire ln_if_47_acc_itm_13_1;
  wire ln_if_46_acc_itm_14_1;
  wire ln_if_45_acc_itm_14_1;
  wire ln_if_44_acc_itm_12_1;
  wire ln_if_43_acc_itm_14_1;
  wire ln_if_42_acc_itm_13_1;
  wire ln_if_41_acc_itm_14_1;
  wire ln_if_40_acc_itm_11_1;
  wire ln_if_39_acc_itm_14_1;
  wire ln_if_38_acc_itm_14_1;
  wire ln_if_37_acc_itm_13_1;
  wire ln_if_36_acc_itm_14_1;
  wire ln_if_35_acc_itm_11_1;
  wire ln_if_34_acc_itm_14_1;
  wire ln_if_33_acc_itm_13_1;
  wire ln_if_32_acc_itm_14_1;
  wire ln_if_31_acc_itm_14_1;
  wire ln_if_30_acc_itm_11_1;
  wire ln_if_29_acc_itm_14_1;
  wire ln_if_28_acc_itm_13_1;
  wire ln_if_27_acc_itm_14_1;
  wire ln_if_26_acc_itm_12_1;
  wire ln_if_25_acc_itm_14_1;
  wire ln_if_24_acc_itm_14_1;
  wire ln_if_23_acc_itm_13_1;
  wire ln_if_22_acc_itm_14_1;
  wire ln_if_21_acc_itm_12_1;
  wire ln_if_20_acc_itm_14_1;
  wire ln_if_19_acc_itm_13_1;
  wire ln_if_18_acc_itm_14_1;
  wire ln_if_17_acc_itm_14_1;
  wire ln_if_16_acc_itm_12_1;
  wire ln_if_15_acc_itm_14_1;
  wire ln_if_14_acc_itm_13_1;
  wire ln_if_13_acc_itm_14_1;
  wire ln_if_12_acc_itm_10_1;
  wire ln_if_11_acc_itm_14_1;
  wire ln_if_10_acc_itm_14_1;
  wire ln_if_9_acc_itm_13_1;
  wire ln_if_8_acc_itm_14_1;
  wire ln_if_4_acc_itm_8_1;
  wire ln_if_5_acc_itm_7_1;
  wire ln_if_3_acc_itm_6_1;
  wire ln_if_2_acc_itm_8_1;
  wire ln_1_if_252_acc_itm_12_1;
  wire ln_1_if_244_acc_itm_14_1;
  wire ln_1_if_245_acc_itm_13_1;
  wire ln_1_if_251_acc_itm_10_1;
  wire ln_1_if_250_acc_itm_12_1;
  wire ln_1_if_249_acc_itm_11_1;
  wire ln_1_if_248_acc_itm_12_1;
  wire ln_1_if_247_acc_itm_9_1;
  wire ln_1_if_246_acc_itm_14_1;
  wire ln_1_if_144_acc_itm_14_1;
  wire ln_1_if_145_acc_itm_13_1;
  wire ln_1_if_243_acc_itm_12_1;
  wire ln_1_if_242_acc_itm_14_1;
  wire ln_1_if_241_acc_itm_13_1;
  wire ln_1_if_240_acc_itm_14_1;
  wire ln_1_if_239_acc_itm_11_1;
  wire ln_1_if_238_acc_itm_14_1;
  wire ln_1_if_237_acc_itm_13_1;
  wire ln_1_if_236_acc_itm_14_1;
  wire ln_1_if_235_acc_itm_12_1;
  wire ln_1_if_234_acc_itm_14_1;
  wire ln_1_if_233_acc_itm_13_1;
  wire ln_1_if_232_acc_itm_14_1;
  wire ln_1_if_231_acc_itm_10_1;
  wire ln_1_if_230_acc_itm_14_1;
  wire ln_1_if_229_acc_itm_13_1;
  wire ln_1_if_228_acc_itm_14_1;
  wire ln_1_if_227_acc_itm_12_1;
  wire ln_1_if_226_acc_itm_14_1;
  wire ln_1_if_225_acc_itm_13_1;
  wire ln_1_if_224_acc_itm_14_1;
  wire ln_1_if_223_acc_itm_11_1;
  wire ln_1_if_222_acc_itm_14_1;
  wire ln_1_if_221_acc_itm_13_1;
  wire ln_1_if_220_acc_itm_14_1;
  wire ln_1_if_219_acc_itm_12_1;
  wire ln_1_if_218_acc_itm_14_1;
  wire ln_1_if_217_acc_itm_13_1;
  wire ln_1_if_216_acc_itm_14_1;
  wire ln_1_if_215_acc_itm_8_1;
  wire ln_1_if_214_acc_itm_14_1;
  wire ln_1_if_213_acc_itm_13_1;
  wire ln_1_if_212_acc_itm_14_1;
  wire ln_1_if_211_acc_itm_12_1;
  wire ln_1_if_210_acc_itm_14_1;
  wire ln_1_if_209_acc_itm_13_1;
  wire ln_1_if_208_acc_itm_14_1;
  wire ln_1_if_207_acc_itm_11_1;
  wire ln_1_if_206_acc_itm_14_1;
  wire ln_1_if_205_acc_itm_13_1;
  wire ln_1_if_204_acc_itm_14_1;
  wire ln_1_if_203_acc_itm_12_1;
  wire ln_1_if_202_acc_itm_14_1;
  wire ln_1_if_201_acc_itm_13_1;
  wire ln_1_if_200_acc_itm_14_1;
  wire ln_1_if_199_acc_itm_10_1;
  wire ln_1_if_198_acc_itm_14_1;
  wire ln_1_if_197_acc_itm_13_1;
  wire ln_1_if_196_acc_itm_14_1;
  wire ln_1_if_195_acc_itm_12_1;
  wire ln_1_if_194_acc_itm_14_1;
  wire ln_1_if_193_acc_itm_13_1;
  wire ln_1_if_192_acc_itm_14_1;
  wire ln_1_if_191_acc_itm_11_1;
  wire ln_1_if_190_acc_itm_14_1;
  wire ln_1_if_189_acc_itm_13_1;
  wire ln_1_if_188_acc_itm_14_1;
  wire ln_1_if_187_acc_itm_12_1;
  wire ln_1_if_186_acc_itm_14_1;
  wire ln_1_if_185_acc_itm_13_1;
  wire ln_1_if_184_acc_itm_14_1;
  wire ln_1_if_183_acc_itm_9_1;
  wire ln_1_if_182_acc_itm_14_1;
  wire ln_1_if_181_acc_itm_13_1;
  wire ln_1_if_180_acc_itm_14_1;
  wire ln_1_if_179_acc_itm_12_1;
  wire ln_1_if_178_acc_itm_14_1;
  wire ln_1_if_177_acc_itm_13_1;
  wire ln_1_if_176_acc_itm_14_1;
  wire ln_1_if_175_acc_itm_11_1;
  wire ln_1_if_174_acc_itm_14_1;
  wire ln_1_if_173_acc_itm_13_1;
  wire ln_1_if_172_acc_itm_14_1;
  wire ln_1_if_171_acc_itm_12_1;
  wire ln_1_if_170_acc_itm_14_1;
  wire ln_1_if_169_acc_itm_13_1;
  wire ln_1_if_168_acc_itm_14_1;
  wire ln_1_if_167_acc_itm_10_1;
  wire ln_1_if_166_acc_itm_14_1;
  wire ln_1_if_165_acc_itm_13_1;
  wire ln_1_if_164_acc_itm_14_1;
  wire ln_1_if_163_acc_itm_12_1;
  wire ln_1_if_162_acc_itm_14_1;
  wire ln_1_if_161_acc_itm_13_1;
  wire ln_1_if_160_acc_itm_14_1;
  wire ln_1_if_159_acc_itm_11_1;
  wire ln_1_if_158_acc_itm_14_1;
  wire ln_1_if_157_acc_itm_13_1;
  wire ln_1_if_156_acc_itm_14_1;
  wire ln_1_if_155_acc_itm_12_1;
  wire ln_1_if_154_acc_itm_14_1;
  wire ln_1_if_153_acc_itm_13_1;
  wire ln_1_if_152_acc_itm_14_1;
  wire ln_1_if_151_acc_itm_7_1;
  wire ln_1_if_150_acc_itm_14_1;
  wire ln_1_if_149_acc_itm_13_1;
  wire ln_1_if_148_acc_itm_14_1;
  wire ln_1_if_147_acc_itm_12_1;
  wire ln_1_if_146_acc_itm_14_1;
  wire ln_1_if_142_acc_itm_14_1;
  wire ln_1_if_143_acc_itm_11_1;
  wire ln_1_if_141_acc_itm_13_1;
  wire ln_1_if_140_acc_itm_14_1;
  wire ln_1_if_52_acc_itm_14_1;
  wire ln_1_if_53_acc_itm_14_1;
  wire ln_1_if_49_acc_itm_12_1;
  wire ln_1_if_50_acc_itm_14_1;
  wire ln_1_if_6_acc_itm_8_1;
  wire ln_1_if_7_acc_itm_5_1;
  wire ln_1_if_139_acc_itm_12_1;
  wire ln_1_if_138_acc_itm_14_1;
  wire ln_1_if_137_acc_itm_13_1;
  wire ln_1_if_136_acc_itm_14_1;
  wire ln_1_if_135_acc_itm_10_1;
  wire ln_1_if_134_acc_itm_14_1;
  wire ln_1_if_133_acc_itm_13_1;
  wire ln_1_if_132_acc_itm_14_1;
  wire ln_1_if_131_acc_itm_12_1;
  wire ln_1_if_130_acc_itm_14_1;
  wire ln_1_if_129_acc_itm_13_1;
  wire ln_1_if_128_acc_itm_14_1;
  wire ln_1_if_127_acc_itm_11_1;
  wire ln_1_if_126_acc_itm_14_1;
  wire ln_1_if_125_acc_itm_13_1;
  wire ln_1_if_124_acc_itm_14_1;
  wire ln_1_if_123_acc_itm_12_1;
  wire ln_1_if_122_acc_itm_14_1;
  wire ln_1_if_121_acc_itm_13_1;
  wire ln_1_if_120_acc_itm_14_1;
  wire ln_1_if_119_acc_itm_9_1;
  wire ln_1_if_118_acc_itm_14_1;
  wire ln_1_if_117_acc_itm_13_1;
  wire ln_1_if_116_acc_itm_14_1;
  wire ln_1_if_115_acc_itm_14_1;
  wire ln_1_if_114_acc_itm_10_1;
  wire ln_1_if_113_acc_itm_14_1;
  wire ln_1_if_112_acc_itm_13_1;
  wire ln_1_if_111_acc_itm_14_1;
  wire ln_1_if_110_acc_itm_12_1;
  wire ln_1_if_109_acc_itm_14_1;
  wire ln_1_if_108_acc_itm_14_1;
  wire ln_1_if_107_acc_itm_13_1;
  wire ln_1_if_106_acc_itm_14_1;
  wire ln_1_if_105_acc_itm_12_1;
  wire ln_1_if_104_acc_itm_14_1;
  wire ln_1_if_103_acc_itm_13_1;
  wire ln_1_if_102_acc_itm_14_1;
  wire ln_1_if_101_acc_itm_14_1;
  wire ln_1_if_100_acc_itm_12_1;
  wire ln_1_if_99_acc_itm_14_1;
  wire ln_1_if_98_acc_itm_13_1;
  wire ln_1_if_97_acc_itm_14_1;
  wire ln_1_if_96_acc_itm_11_1;
  wire ln_1_if_95_acc_itm_14_1;
  wire ln_1_if_94_acc_itm_14_1;
  wire ln_1_if_93_acc_itm_13_1;
  wire ln_1_if_92_acc_itm_14_1;
  wire ln_1_if_91_acc_itm_11_1;
  wire ln_1_if_90_acc_itm_14_1;
  wire ln_1_if_89_acc_itm_13_1;
  wire ln_1_if_88_acc_itm_14_1;
  wire ln_1_if_87_acc_itm_14_1;
  wire ln_1_if_86_acc_itm_11_1;
  wire ln_1_if_85_acc_itm_14_1;
  wire ln_1_if_84_acc_itm_13_1;
  wire ln_1_if_83_acc_itm_14_1;
  wire ln_1_if_82_acc_itm_12_1;
  wire ln_1_if_81_acc_itm_14_1;
  wire ln_1_if_80_acc_itm_14_1;
  wire ln_1_if_79_acc_itm_13_1;
  wire ln_1_if_78_acc_itm_14_1;
  wire ln_1_if_77_acc_itm_12_1;
  wire ln_1_if_76_acc_itm_14_1;
  wire ln_1_if_75_acc_itm_13_1;
  wire ln_1_if_74_acc_itm_14_1;
  wire ln_1_if_73_acc_itm_14_1;
  wire ln_1_if_72_acc_itm_12_1;
  wire ln_1_if_71_acc_itm_14_1;
  wire ln_1_if_70_acc_itm_13_1;
  wire ln_1_if_69_acc_itm_14_1;
  wire ln_1_if_68_acc_itm_8_1;
  wire ln_1_if_67_acc_itm_14_1;
  wire ln_1_if_66_acc_itm_14_1;
  wire ln_1_if_65_acc_itm_13_1;
  wire ln_1_if_64_acc_itm_14_1;
  wire ln_1_if_63_acc_itm_10_1;
  wire ln_1_if_62_acc_itm_14_1;
  wire ln_1_if_61_acc_itm_13_1;
  wire ln_1_if_60_acc_itm_14_1;
  wire ln_1_if_59_acc_itm_14_1;
  wire ln_1_if_58_acc_itm_9_1;
  wire ln_1_if_57_acc_itm_14_1;
  wire ln_1_if_56_acc_itm_13_1;
  wire ln_1_if_55_acc_itm_14_1;
  wire ln_1_if_54_acc_itm_12_1;
  wire ln_1_if_51_acc_itm_13_1;
  wire ln_1_if_48_acc_itm_14_1;
  wire ln_1_if_47_acc_itm_13_1;
  wire ln_1_if_46_acc_itm_14_1;
  wire ln_1_if_45_acc_itm_14_1;
  wire ln_1_if_44_acc_itm_12_1;
  wire ln_1_if_43_acc_itm_14_1;
  wire ln_1_if_42_acc_itm_13_1;
  wire ln_1_if_41_acc_itm_14_1;
  wire ln_1_if_40_acc_itm_11_1;
  wire ln_1_if_39_acc_itm_14_1;
  wire ln_1_if_38_acc_itm_14_1;
  wire ln_1_if_37_acc_itm_13_1;
  wire ln_1_if_36_acc_itm_14_1;
  wire ln_1_if_35_acc_itm_11_1;
  wire ln_1_if_34_acc_itm_14_1;
  wire ln_1_if_33_acc_itm_13_1;
  wire ln_1_if_32_acc_itm_14_1;
  wire ln_1_if_31_acc_itm_14_1;
  wire ln_1_if_30_acc_itm_11_1;
  wire ln_1_if_29_acc_itm_14_1;
  wire ln_1_if_28_acc_itm_13_1;
  wire ln_1_if_27_acc_itm_14_1;
  wire ln_1_if_26_acc_itm_12_1;
  wire ln_1_if_25_acc_itm_14_1;
  wire ln_1_if_24_acc_itm_14_1;
  wire ln_1_if_23_acc_itm_13_1;
  wire ln_1_if_22_acc_itm_14_1;
  wire ln_1_if_21_acc_itm_12_1;
  wire ln_1_if_20_acc_itm_14_1;
  wire ln_1_if_19_acc_itm_13_1;
  wire ln_1_if_18_acc_itm_14_1;
  wire ln_1_if_17_acc_itm_14_1;
  wire ln_1_if_16_acc_itm_12_1;
  wire ln_1_if_15_acc_itm_14_1;
  wire ln_1_if_14_acc_itm_13_1;
  wire ln_1_if_13_acc_itm_14_1;
  wire ln_1_if_12_acc_itm_10_1;
  wire ln_1_if_11_acc_itm_14_1;
  wire ln_1_if_10_acc_itm_14_1;
  wire ln_1_if_9_acc_itm_13_1;
  wire ln_1_if_8_acc_itm_14_1;
  wire ln_1_if_4_acc_itm_8_1;
  wire ln_1_if_5_acc_itm_7_1;
  wire ln_1_if_3_acc_itm_6_1;
  wire ln_1_if_2_acc_itm_8_1;
  reg [1:0] P1_0_1_23_10_sva_rsp_0;
  reg [11:0] P1_0_1_23_10_sva_rsp_1;
  wire mux_1772_ssc;
  wire or_98_ssc;
  wire [1:0] P1_0_1_23_10_sva_dfm_1_mx0_13_12;
  wire [11:0] P1_0_1_23_10_sva_dfm_1_mx0_11_0;
  wire nand_53_ssc;
  wire and_76_ssc;
  wire and_8_ssc;
  wire [1:0] P1_0_1_23_10_sva_dfm_3_13_12;
  wire [11:0] P1_0_1_23_10_sva_dfm_3_11_0;

  wire[13:0] if_4_aelse_acc_nl;
  wire[14:0] nl_if_4_aelse_acc_nl;
  wire or_40_nl;
  wire if_4_for_if_4_for_if_4_for_not_1_nl;
  wire and_275_nl;
  wire if_4_for_if_4_for_if_4_for_not_2_nl;
  wire and_277_nl;
  wire[13:0] if_4_for_1_and_52_nl;
  wire if_4_for_1_if_4_for_1_nand_1_nl;
  wire mux_1430_nl;
  wire mux_1429_nl;
  wire nand_91_nl;
  wire mux_1428_nl;
  wire mux_1427_nl;
  wire mux_1420_nl;
  wire mux_1419_nl;
  wire[13:0] if_4_for_1_and_44_nl;
  wire if_4_for_1_if_4_for_1_nand_14_nl;
  wire[13:0] if_4_for_1_and_53_nl;
  wire if_4_for_1_if_4_for_1_nand_3_nl;
  wire mux_1453_nl;
  wire mux_1452_nl;
  wire nand_93_nl;
  wire mux_1451_nl;
  wire mux_1450_nl;
  wire mux_1445_nl;
  wire mux_1444_nl;
  wire[13:0] if_4_for_1_and_45_nl;
  wire if_4_for_1_if_4_for_1_nand_12_nl;
  wire mux_1466_nl;
  wire mux_1465_nl;
  wire mux_1464_nl;
  wire nand_70_nl;
  wire mux_1463_nl;
  wire mux_1462_nl;
  wire mux_1461_nl;
  wire mux_1460_nl;
  wire mux_1459_nl;
  wire[13:0] if_4_for_1_and_54_nl;
  wire if_4_for_1_if_4_for_1_nand_5_nl;
  wire mux_1484_nl;
  wire mux_1483_nl;
  wire nand_95_nl;
  wire mux_1482_nl;
  wire mux_1481_nl;
  wire mux_1477_nl;
  wire mux_1476_nl;
  wire[13:0] if_4_for_1_and_46_nl;
  wire if_4_for_1_if_4_for_1_nand_10_nl;
  wire mux_1510_nl;
  wire mux_1509_nl;
  wire nand_96_nl;
  wire mux_1508_nl;
  wire mux_1507_nl;
  wire mux_1501_nl;
  wire mux_1500_nl;
  wire mux_1498_nl;
  wire mux_1497_nl;
  wire mux_1489_nl;
  wire mux_1488_nl;
  wire[13:0] if_4_for_1_and_55_nl;
  wire if_4_for_1_if_4_for_1_nand_7_nl;
  wire mux_1540_nl;
  wire mux_1539_nl;
  wire nand_98_nl;
  wire mux_1538_nl;
  wire mux_1537_nl;
  wire mux_1523_nl;
  wire mux_1522_nl;
  wire[13:0] if_4_for_1_and_47_nl;
  wire if_4_for_1_if_4_for_1_nand_8_nl;
  wire mux_1568_nl;
  wire mux_1567_nl;
  wire nand_99_nl;
  wire mux_1566_nl;
  wire mux_1565_nl;
  wire mux_1555_nl;
  wire mux_1554_nl;
  wire mux_1552_nl;
  wire mux_1551_nl;
  wire mux_1542_nl;
  wire[13:0] if_4_for_1_and_56_nl;
  wire if_4_for_1_if_4_for_1_nand_9_nl;
  wire mux_1596_nl;
  wire mux_1595_nl;
  wire or_434_nl;
  wire mux_1594_nl;
  wire mux_1593_nl;
  wire mux_1583_nl;
  wire mux_1582_nl;
  wire mux_1580_nl;
  wire mux_1579_nl;
  wire mux_1570_nl;
  wire[13:0] if_4_for_1_and_48_nl;
  wire if_4_for_1_if_4_for_1_nand_6_nl;
  wire mux_1625_nl;
  wire mux_1624_nl;
  wire nand_102_nl;
  wire mux_1623_nl;
  wire mux_1622_nl;
  wire mux_1609_nl;
  wire mux_1608_nl;
  wire[13:0] if_4_for_1_and_57_nl;
  wire if_4_for_1_if_4_for_1_nand_11_nl;
  wire mux_1656_nl;
  wire mux_1655_nl;
  wire or_469_nl;
  wire mux_1654_nl;
  wire mux_1653_nl;
  wire mux_1645_nl;
  wire mux_1644_nl;
  wire mux_1641_nl;
  wire mux_1640_nl;
  wire mux_1631_nl;
  wire mux_1628_nl;
  wire[13:0] if_4_for_1_and_49_nl;
  wire if_4_for_1_if_4_for_1_nand_4_nl;
  wire mux_1673_nl;
  wire mux_1672_nl;
  wire nand_105_nl;
  wire mux_1671_nl;
  wire mux_1670_nl;
  wire mux_1665_nl;
  wire mux_1664_nl;
  wire[13:0] if_4_for_1_and_58_nl;
  wire if_4_for_1_if_4_for_1_nand_13_nl;
  wire mux_1695_nl;
  wire mux_1694_nl;
  wire or_498_nl;
  wire mux_1693_nl;
  wire mux_1692_nl;
  wire mux_1681_nl;
  wire mux_1680_nl;
  wire[13:0] if_4_for_1_and_50_nl;
  wire if_4_for_1_if_4_for_1_nand_2_nl;
  wire mux_1718_nl;
  wire mux_1717_nl;
  wire nand_108_nl;
  wire mux_1716_nl;
  wire mux_1715_nl;
  wire mux_1710_nl;
  wire mux_1709_nl;
  wire[13:0] if_4_for_1_and_59_nl;
  wire if_4_for_1_if_4_for_1_nand_15_nl;
  wire mux_1726_nl;
  wire and_283_nl;
  wire mux_1725_nl;
  wire mux_1724_nl;
  wire and_285_nl;
  wire and_286_nl;
  wire and_258_nl;
  wire[13:0] if_4_for_1_and_51_nl;
  wire if_4_for_1_if_4_for_1_nand_nl;
  wire mux_1750_nl;
  wire mux_1749_nl;
  wire nand_109_nl;
  wire mux_1748_nl;
  wire mux_1747_nl;
  wire mux_1740_nl;
  wire mux_1739_nl;
  wire nor_67_nl;
  wire mux_1769_nl;
  wire mux_1768_nl;
  wire mux_1767_nl;
  wire or_545_nl;
  wire mux_1766_nl;
  wire mux_1765_nl;
  wire mux_1764_nl;
  wire mux_1763_nl;
  wire mux_1762_nl;
  wire mux_1761_nl;
  wire mux_1760_nl;
  wire mux_1759_nl;
  wire mux_1758_nl;
  wire nor_68_nl;
  wire mux_1791_nl;
  wire mux_1790_nl;
  wire mux_1789_nl;
  wire or_564_nl;
  wire mux_1788_nl;
  wire mux_1787_nl;
  wire mux_1786_nl;
  wire mux_1785_nl;
  wire mux_1784_nl;
  wire nand_110_nl;
  wire if_4_for_if_4_for_nand_4_nl;
  wire nor_69_nl;
  wire mux_1809_nl;
  wire mux_1808_nl;
  wire nand_83_nl;
  wire mux_1807_nl;
  wire mux_1806_nl;
  wire mux_1805_nl;
  wire mux_1804_nl;
  wire mux_1803_nl;
  wire mux_1802_nl;
  wire mux_1801_nl;
  wire mux_1797_nl;
  wire mux_1796_nl;
  wire mux_1795_nl;
  wire mux_1794_nl;
  wire nor_70_nl;
  wire mux_1826_nl;
  wire mux_1825_nl;
  wire or_581_nl;
  wire mux_1824_nl;
  wire mux_1823_nl;
  wire mux_1821_nl;
  wire mux_1820_nl;
  wire mux_1819_nl;
  wire mux_1818_nl;
  wire mux_1817_nl;
  wire mux_1815_nl;
  wire mux_1814_nl;
  wire mux_1813_nl;
  wire mux_1812_nl;
  wire if_4_for_if_4_for_nand_2_nl;
  wire nor_71_nl;
  wire mux_1845_nl;
  wire mux_1844_nl;
  wire mux_1843_nl;
  wire or_608_nl;
  wire mux_1842_nl;
  wire mux_1841_nl;
  wire mux_1840_nl;
  wire mux_1839_nl;
  wire mux_1838_nl;
  wire or_583_nl;
  wire nor_72_nl;
  wire mux_1854_nl;
  wire and_293_nl;
  wire mux_1853_nl;
  wire and_263_nl;
  wire mux_1852_nl;
  wire if_4_for_if_4_for_nand_nl;
  wire nor_73_nl;
  wire mux_1874_nl;
  wire mux_1873_nl;
  wire mux_1872_nl;
  wire nand_88_nl;
  wire mux_1871_nl;
  wire mux_1870_nl;
  wire mux_1869_nl;
  wire mux_1868_nl;
  wire mux_1867_nl;
  wire mux_1866_nl;
  wire mux_1865_nl;
  wire mux_1864_nl;
  wire mux_1863_nl;
  wire not_402_nl;
  wire mux_1306_nl;
  wire nor_51_nl;
  wire if_4_for_if_4_for_or_4_nl;
  wire[15:0] if_4_acc_1_nl;
  wire[16:0] nl_if_4_acc_1_nl;
  wire[11:0] ln_if_253_acc_nl;
  wire[12:0] nl_ln_if_253_acc_nl;
  wire[14:0] operator_24_14_false_AC_TRN_AC_WRAP_acc_nl;
  wire[15:0] nl_operator_24_14_false_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] ln_1_if_253_acc_nl;
  wire[12:0] nl_ln_1_if_253_acc_nl;
  wire[23:0] if_4_for_if_acc_nl;
  wire[24:0] nl_if_4_for_if_acc_nl;
  wire[24:0] if_4_for_if_if_4_for_if_mul_nl;
  wire signed [29:0] nl_if_4_for_if_if_4_for_if_mul_nl;
  wire ln_ln_ln_and_4_nl;
  wire ln_ln_ln_or_20_nl;
  wire ln_ln_ln_or_21_nl;
  wire ln_ln_ln_and_5_nl;
  wire ln_ln_ln_or_24_nl;
  wire ln_ln_ln_or_26_nl;
  wire ln_ln_ln_or_27_nl;
  wire ln_ln_ln_and_6_nl;
  wire ln_ln_ln_or_30_nl;
  wire ln_ln_ln_and_7_nl;
  wire ln_ln_ln_or_32_nl;
  wire ln_ln_ln_or_34_nl;
  wire ln_ln_ln_or_36_nl;
  wire ln_ln_ln_or_37_nl;
  wire[23:0] if_4_for_1_if_acc_nl;
  wire[24:0] nl_if_4_for_1_if_acc_nl;
  wire[24:0] if_4_for_1_if_if_4_for_1_if_mul_nl;
  wire signed [29:0] nl_if_4_for_1_if_if_4_for_1_if_mul_nl;
  wire ln_1_ln_1_ln_1_and_4_nl;
  wire ln_1_ln_1_ln_1_or_20_nl;
  wire ln_1_ln_1_ln_1_or_21_nl;
  wire ln_1_ln_1_ln_1_and_5_nl;
  wire ln_1_ln_1_ln_1_or_24_nl;
  wire ln_1_ln_1_ln_1_or_26_nl;
  wire ln_1_ln_1_ln_1_or_27_nl;
  wire ln_1_ln_1_ln_1_and_6_nl;
  wire ln_1_ln_1_ln_1_or_30_nl;
  wire ln_1_ln_1_ln_1_and_7_nl;
  wire ln_1_ln_1_ln_1_or_32_nl;
  wire ln_1_ln_1_ln_1_or_34_nl;
  wire ln_1_ln_1_ln_1_or_36_nl;
  wire ln_1_ln_1_ln_1_or_37_nl;
  wire[14:0] operator_24_14_false_AC_TRN_AC_WRAP_1_acc_nl;
  wire[15:0] nl_operator_24_14_false_AC_TRN_AC_WRAP_1_acc_nl;
  wire or_49_nl;
  wire or_55_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_operator_24_14_false_AC_TRN_AC_WRAP_operator_24_14_false_AC_TRN_AC_WRAP_mux_nl;
  wire or_58_nl;
  wire or_61_nl;
  wire or_65_nl;
  wire or_68_nl;
  wire or_70_nl;
  wire or_72_nl;
  wire or_76_nl;
  wire or_79_nl;
  wire or_81_nl;
  wire or_83_nl;
  wire or_87_nl;
  wire or_90_nl;
  wire or_92_nl;
  wire or_94_nl;
  wire or_102_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_nl;
  wire or_104_nl;
  wire or_106_nl;
  wire or_109_nl;
  wire or_112_nl;
  wire or_114_nl;
  wire or_116_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_6_operator_24_14_false_AC_TRN_AC_WRAP_6_operator_24_14_false_AC_TRN_AC_WRAP_6_mux_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_mux_3_nl;
  wire or_135_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_mux_7_nl;
  wire or_142_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_mux_11_nl;
  wire or_153_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_mux_15_nl;
  wire or_159_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_mux_19_nl;
  wire or_169_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_mux_23_nl;
  wire or_177_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_mux_27_nl;
  wire or_184_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_mux_31_nl;
  wire or_192_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_mux_1_nl;
  wire or_129_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_mux_5_nl;
  wire or_140_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_mux_9_nl;
  wire or_151_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_mux_13_nl;
  wire or_157_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_mux_17_nl;
  wire or_162_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_mux_21_nl;
  wire or_171_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_mux_25_nl;
  wire or_179_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_mux_29_nl;
  wire or_189_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_3_operator_24_14_false_AC_TRN_AC_WRAP_3_operator_24_14_false_AC_TRN_AC_WRAP_3_operator_24_14_false_AC_TRN_AC_WRAP_3_mux1h_nl;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_12_nl;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_or_nl;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_or_1_nl;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_35_nl;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_37_nl;
  wire operator_24_14_false_AC_TRN_AC_WRAP_3_and_27_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_2_operator_24_14_false_AC_TRN_AC_WRAP_2_operator_24_14_false_AC_TRN_AC_WRAP_2_operator_24_14_false_AC_TRN_AC_WRAP_2_mux1h_nl;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_or_nl;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_20_nl;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_21_nl;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_22_nl;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_23_nl;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_25_nl;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_26_nl;
  wire operator_24_14_false_AC_TRN_AC_WRAP_2_and_27_nl;
  wire or_195_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_5_operator_24_14_false_AC_TRN_AC_WRAP_5_operator_24_14_false_AC_TRN_AC_WRAP_5_mux_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_mux_3_nl;
  wire or_202_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_mux_7_nl;
  wire or_206_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_mux_11_nl;
  wire or_216_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_mux_15_nl;
  wire or_230_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_mux_19_nl;
  wire or_246_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_mux_23_nl;
  wire or_256_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_mux_27_nl;
  wire or_264_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_mux_31_nl;
  wire or_269_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_mux_29_nl;
  wire or_266_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_mux_25_nl;
  wire or_260_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_mux_21_nl;
  wire or_252_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_mux_17_nl;
  wire or_237_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_mux_13_nl;
  wire or_224_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_mux_9_nl;
  wire or_213_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_mux_5_nl;
  wire or_204_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_mux_1_nl;
  wire or_197_nl;
  wire or_200_nl;
  wire or_203_nl;
  wire mux_1354_nl;
  wire or_205_nl;
  wire mux_1355_nl;
  wire or_211_nl;
  wire mux_1363_nl;
  wire mux_1359_nl;
  wire or_214_nl;
  wire mux_1365_nl;
  wire mux_1364_nl;
  wire or_221_nl;
  wire or_219_nl;
  wire or_223_nl;
  wire mux_1369_nl;
  wire and_183_nl;
  wire or_229_nl;
  wire mux_1373_nl;
  wire mux_1370_nl;
  wire or_225_nl;
  wire nand_45_nl;
  wire mux_1377_nl;
  wire mux_1374_nl;
  wire nor_64_nl;
  wire or_244_nl;
  wire mux_1381_nl;
  wire or_295_nl;
  wire mux_1384_nl;
  wire or_249_nl;
  wire mux_1387_nl;
  wire or_293_nl;
  wire or_258_nl;
  wire mux_1388_nl;
  wire or_262_nl;
  wire mux_1389_nl;
  wire or_265_nl;
  wire mux_1390_nl;
  wire nand_9_nl;
  wire or_268_nl;
  wire mux_1391_nl;
  wire or_267_nl;
  wire[13:0] operator_24_14_false_AC_TRN_AC_WRAP_4_operator_24_14_false_AC_TRN_AC_WRAP_4_operator_24_14_false_AC_TRN_AC_WRAP_4_mux_nl;
  wire nor_66_nl;
  wire if_4_for_if_4_for_if_4_for_not_3_nl;
  wire nand_55_nl;
  wire and_78_nl;
  wire and_10_nl;
  wire nand_57_nl;
  wire and_80_nl;
  wire and_12_nl;
  wire nand_59_nl;
  wire and_82_nl;
  wire and_14_nl;
  wire nand_61_nl;
  wire and_84_nl;
  wire and_16_nl;
  wire nand_63_nl;
  wire and_86_nl;
  wire and_18_nl;
  wire nand_65_nl;
  wire and_88_nl;
  wire and_20_nl;
  wire nand_67_nl;
  wire and_90_nl;
  wire and_22_nl;
  wire if_4_for_if_4_for_if_4_for_not_20_nl;
  wire and_200_nl;
  wire and_201_nl;
  wire and_24_nl;
  wire mux_1322_nl;
  wire and_202_nl;
  wire and_203_nl;
  wire and_26_nl;
  wire mux_1331_nl;
  wire mux_1330_nl;
  wire and_204_nl;
  wire and_205_nl;
  wire and_28_nl;
  wire mux_1337_nl;
  wire and_206_nl;
  wire and_207_nl;
  wire and_30_nl;
  wire mux_1341_nl;
  wire or_166_nl;
  wire mux_1340_nl;
  wire or_165_nl;
  wire and_208_nl;
  wire and_209_nl;
  wire and_32_nl;
  wire mux_1345_nl;
  wire or_176_nl;
  wire or_175_nl;
  wire or_173_nl;
  wire and_210_nl;
  wire and_211_nl;
  wire and_34_nl;
  wire mux_1350_nl;
  wire nand_4_nl;
  wire mux_1349_nl;
  wire or_182_nl;
  wire and_212_nl;
  wire and_213_nl;
  wire and_36_nl;
  wire nand_5_nl;
  wire mux_1352_nl;
  wire or_191_nl;
  wire and_214_nl;
  wire and_215_nl;
  wire and_38_nl;
  wire or_122_nl;
  wire mux_1312_nl;
  wire or_120_nl;
  wire and_216_nl;
  wire and_217_nl;
  wire and_40_nl;
  wire mux_1319_nl;
  wire nor_61_nl;
  wire mux_1318_nl;
  wire nor_62_nl;
  wire and_218_nl;
  wire and_219_nl;
  wire and_42_nl;
  wire or_149_nl;
  wire mux_1324_nl;
  wire or_147_nl;
  wire or_145_nl;
  wire and_220_nl;
  wire and_221_nl;
  wire and_44_nl;
  wire mux_1334_nl;
  wire and_197_nl;
  wire mux_1333_nl;
  wire and_198_nl;
  wire and_222_nl;
  wire and_223_nl;
  wire and_46_nl;
  wire mux_1338_nl;
  wire and_224_nl;
  wire and_225_nl;
  wire and_48_nl;
  wire mux_1343_nl;
  wire mux_1342_nl;
  wire and_226_nl;
  wire and_227_nl;
  wire and_50_nl;
  wire mux_1347_nl;
  wire and_228_nl;
  wire and_229_nl;
  wire and_52_nl;
  wire and_230_nl;
  wire and_231_nl;
  wire and_54_nl;
  wire or_288_nl;
  wire[12:0] ln_if_252_acc_nl;
  wire[13:0] nl_ln_if_252_acc_nl;
  wire[14:0] ln_if_244_acc_nl;
  wire[15:0] nl_ln_if_244_acc_nl;
  wire[13:0] ln_if_245_acc_nl;
  wire[14:0] nl_ln_if_245_acc_nl;
  wire[10:0] ln_if_251_acc_nl;
  wire[11:0] nl_ln_if_251_acc_nl;
  wire[12:0] ln_if_250_acc_nl;
  wire[13:0] nl_ln_if_250_acc_nl;
  wire[11:0] ln_if_249_acc_nl;
  wire[12:0] nl_ln_if_249_acc_nl;
  wire[12:0] ln_if_248_acc_nl;
  wire[13:0] nl_ln_if_248_acc_nl;
  wire[9:0] ln_if_247_acc_nl;
  wire[10:0] nl_ln_if_247_acc_nl;
  wire[14:0] ln_if_246_acc_nl;
  wire[15:0] nl_ln_if_246_acc_nl;
  wire[7:0] ln_if_1_acc_nl;
  wire[8:0] nl_ln_if_1_acc_nl;
  wire[14:0] ln_if_144_acc_nl;
  wire[15:0] nl_ln_if_144_acc_nl;
  wire[13:0] ln_if_145_acc_nl;
  wire[14:0] nl_ln_if_145_acc_nl;
  wire[12:0] ln_if_243_acc_nl;
  wire[13:0] nl_ln_if_243_acc_nl;
  wire[14:0] ln_if_242_acc_nl;
  wire[15:0] nl_ln_if_242_acc_nl;
  wire[13:0] ln_if_241_acc_nl;
  wire[14:0] nl_ln_if_241_acc_nl;
  wire[14:0] ln_if_240_acc_nl;
  wire[15:0] nl_ln_if_240_acc_nl;
  wire[11:0] ln_if_239_acc_nl;
  wire[12:0] nl_ln_if_239_acc_nl;
  wire[14:0] ln_if_238_acc_nl;
  wire[15:0] nl_ln_if_238_acc_nl;
  wire[13:0] ln_if_237_acc_nl;
  wire[14:0] nl_ln_if_237_acc_nl;
  wire[14:0] ln_if_236_acc_nl;
  wire[15:0] nl_ln_if_236_acc_nl;
  wire[12:0] ln_if_235_acc_nl;
  wire[13:0] nl_ln_if_235_acc_nl;
  wire[14:0] ln_if_234_acc_nl;
  wire[15:0] nl_ln_if_234_acc_nl;
  wire[13:0] ln_if_233_acc_nl;
  wire[14:0] nl_ln_if_233_acc_nl;
  wire[14:0] ln_if_232_acc_nl;
  wire[15:0] nl_ln_if_232_acc_nl;
  wire[10:0] ln_if_231_acc_nl;
  wire[11:0] nl_ln_if_231_acc_nl;
  wire[14:0] ln_if_230_acc_nl;
  wire[15:0] nl_ln_if_230_acc_nl;
  wire[13:0] ln_if_229_acc_nl;
  wire[14:0] nl_ln_if_229_acc_nl;
  wire[14:0] ln_if_228_acc_nl;
  wire[15:0] nl_ln_if_228_acc_nl;
  wire[12:0] ln_if_227_acc_nl;
  wire[13:0] nl_ln_if_227_acc_nl;
  wire[14:0] ln_if_226_acc_nl;
  wire[15:0] nl_ln_if_226_acc_nl;
  wire[13:0] ln_if_225_acc_nl;
  wire[14:0] nl_ln_if_225_acc_nl;
  wire[14:0] ln_if_224_acc_nl;
  wire[15:0] nl_ln_if_224_acc_nl;
  wire[11:0] ln_if_223_acc_nl;
  wire[12:0] nl_ln_if_223_acc_nl;
  wire[14:0] ln_if_222_acc_nl;
  wire[15:0] nl_ln_if_222_acc_nl;
  wire[13:0] ln_if_221_acc_nl;
  wire[14:0] nl_ln_if_221_acc_nl;
  wire[14:0] ln_if_220_acc_nl;
  wire[15:0] nl_ln_if_220_acc_nl;
  wire[12:0] ln_if_219_acc_nl;
  wire[13:0] nl_ln_if_219_acc_nl;
  wire[14:0] ln_if_218_acc_nl;
  wire[15:0] nl_ln_if_218_acc_nl;
  wire[13:0] ln_if_217_acc_nl;
  wire[14:0] nl_ln_if_217_acc_nl;
  wire[14:0] ln_if_216_acc_nl;
  wire[15:0] nl_ln_if_216_acc_nl;
  wire[8:0] ln_if_215_acc_nl;
  wire[9:0] nl_ln_if_215_acc_nl;
  wire[14:0] ln_if_214_acc_nl;
  wire[15:0] nl_ln_if_214_acc_nl;
  wire[13:0] ln_if_213_acc_nl;
  wire[14:0] nl_ln_if_213_acc_nl;
  wire[14:0] ln_if_212_acc_nl;
  wire[15:0] nl_ln_if_212_acc_nl;
  wire[12:0] ln_if_211_acc_nl;
  wire[13:0] nl_ln_if_211_acc_nl;
  wire[14:0] ln_if_210_acc_nl;
  wire[15:0] nl_ln_if_210_acc_nl;
  wire[13:0] ln_if_209_acc_nl;
  wire[14:0] nl_ln_if_209_acc_nl;
  wire[14:0] ln_if_208_acc_nl;
  wire[15:0] nl_ln_if_208_acc_nl;
  wire[11:0] ln_if_207_acc_nl;
  wire[12:0] nl_ln_if_207_acc_nl;
  wire[14:0] ln_if_206_acc_nl;
  wire[15:0] nl_ln_if_206_acc_nl;
  wire[13:0] ln_if_205_acc_nl;
  wire[14:0] nl_ln_if_205_acc_nl;
  wire[14:0] ln_if_204_acc_nl;
  wire[15:0] nl_ln_if_204_acc_nl;
  wire[12:0] ln_if_203_acc_nl;
  wire[13:0] nl_ln_if_203_acc_nl;
  wire[14:0] ln_if_202_acc_nl;
  wire[15:0] nl_ln_if_202_acc_nl;
  wire[13:0] ln_if_201_acc_nl;
  wire[14:0] nl_ln_if_201_acc_nl;
  wire[14:0] ln_if_200_acc_nl;
  wire[15:0] nl_ln_if_200_acc_nl;
  wire[10:0] ln_if_199_acc_nl;
  wire[11:0] nl_ln_if_199_acc_nl;
  wire[14:0] ln_if_198_acc_nl;
  wire[15:0] nl_ln_if_198_acc_nl;
  wire[13:0] ln_if_197_acc_nl;
  wire[14:0] nl_ln_if_197_acc_nl;
  wire[14:0] ln_if_196_acc_nl;
  wire[15:0] nl_ln_if_196_acc_nl;
  wire[12:0] ln_if_195_acc_nl;
  wire[13:0] nl_ln_if_195_acc_nl;
  wire[14:0] ln_if_194_acc_nl;
  wire[15:0] nl_ln_if_194_acc_nl;
  wire[13:0] ln_if_193_acc_nl;
  wire[14:0] nl_ln_if_193_acc_nl;
  wire[14:0] ln_if_192_acc_nl;
  wire[15:0] nl_ln_if_192_acc_nl;
  wire[11:0] ln_if_191_acc_nl;
  wire[12:0] nl_ln_if_191_acc_nl;
  wire[14:0] ln_if_190_acc_nl;
  wire[15:0] nl_ln_if_190_acc_nl;
  wire[13:0] ln_if_189_acc_nl;
  wire[14:0] nl_ln_if_189_acc_nl;
  wire[14:0] ln_if_188_acc_nl;
  wire[15:0] nl_ln_if_188_acc_nl;
  wire[12:0] ln_if_187_acc_nl;
  wire[13:0] nl_ln_if_187_acc_nl;
  wire[14:0] ln_if_186_acc_nl;
  wire[15:0] nl_ln_if_186_acc_nl;
  wire[13:0] ln_if_185_acc_nl;
  wire[14:0] nl_ln_if_185_acc_nl;
  wire[14:0] ln_if_184_acc_nl;
  wire[15:0] nl_ln_if_184_acc_nl;
  wire[9:0] ln_if_183_acc_nl;
  wire[10:0] nl_ln_if_183_acc_nl;
  wire[14:0] ln_if_182_acc_nl;
  wire[15:0] nl_ln_if_182_acc_nl;
  wire[13:0] ln_if_181_acc_nl;
  wire[14:0] nl_ln_if_181_acc_nl;
  wire[14:0] ln_if_180_acc_nl;
  wire[15:0] nl_ln_if_180_acc_nl;
  wire[12:0] ln_if_179_acc_nl;
  wire[13:0] nl_ln_if_179_acc_nl;
  wire[14:0] ln_if_178_acc_nl;
  wire[15:0] nl_ln_if_178_acc_nl;
  wire[13:0] ln_if_177_acc_nl;
  wire[14:0] nl_ln_if_177_acc_nl;
  wire[14:0] ln_if_176_acc_nl;
  wire[15:0] nl_ln_if_176_acc_nl;
  wire[11:0] ln_if_175_acc_nl;
  wire[12:0] nl_ln_if_175_acc_nl;
  wire[14:0] ln_if_174_acc_nl;
  wire[15:0] nl_ln_if_174_acc_nl;
  wire[13:0] ln_if_173_acc_nl;
  wire[14:0] nl_ln_if_173_acc_nl;
  wire[14:0] ln_if_172_acc_nl;
  wire[15:0] nl_ln_if_172_acc_nl;
  wire[12:0] ln_if_171_acc_nl;
  wire[13:0] nl_ln_if_171_acc_nl;
  wire[14:0] ln_if_170_acc_nl;
  wire[15:0] nl_ln_if_170_acc_nl;
  wire[13:0] ln_if_169_acc_nl;
  wire[14:0] nl_ln_if_169_acc_nl;
  wire[14:0] ln_if_168_acc_nl;
  wire[15:0] nl_ln_if_168_acc_nl;
  wire[10:0] ln_if_167_acc_nl;
  wire[11:0] nl_ln_if_167_acc_nl;
  wire[14:0] ln_if_166_acc_nl;
  wire[15:0] nl_ln_if_166_acc_nl;
  wire[13:0] ln_if_165_acc_nl;
  wire[14:0] nl_ln_if_165_acc_nl;
  wire[14:0] ln_if_164_acc_nl;
  wire[15:0] nl_ln_if_164_acc_nl;
  wire[12:0] ln_if_163_acc_nl;
  wire[13:0] nl_ln_if_163_acc_nl;
  wire[14:0] ln_if_162_acc_nl;
  wire[15:0] nl_ln_if_162_acc_nl;
  wire[13:0] ln_if_161_acc_nl;
  wire[14:0] nl_ln_if_161_acc_nl;
  wire[14:0] ln_if_160_acc_nl;
  wire[15:0] nl_ln_if_160_acc_nl;
  wire[11:0] ln_if_159_acc_nl;
  wire[12:0] nl_ln_if_159_acc_nl;
  wire[14:0] ln_if_158_acc_nl;
  wire[15:0] nl_ln_if_158_acc_nl;
  wire[13:0] ln_if_157_acc_nl;
  wire[14:0] nl_ln_if_157_acc_nl;
  wire[14:0] ln_if_156_acc_nl;
  wire[15:0] nl_ln_if_156_acc_nl;
  wire[12:0] ln_if_155_acc_nl;
  wire[13:0] nl_ln_if_155_acc_nl;
  wire[14:0] ln_if_154_acc_nl;
  wire[15:0] nl_ln_if_154_acc_nl;
  wire[13:0] ln_if_153_acc_nl;
  wire[14:0] nl_ln_if_153_acc_nl;
  wire[14:0] ln_if_152_acc_nl;
  wire[15:0] nl_ln_if_152_acc_nl;
  wire[7:0] ln_if_151_acc_nl;
  wire[8:0] nl_ln_if_151_acc_nl;
  wire[14:0] ln_if_150_acc_nl;
  wire[15:0] nl_ln_if_150_acc_nl;
  wire[13:0] ln_if_149_acc_nl;
  wire[14:0] nl_ln_if_149_acc_nl;
  wire[14:0] ln_if_148_acc_nl;
  wire[15:0] nl_ln_if_148_acc_nl;
  wire[12:0] ln_if_147_acc_nl;
  wire[13:0] nl_ln_if_147_acc_nl;
  wire[14:0] ln_if_146_acc_nl;
  wire[15:0] nl_ln_if_146_acc_nl;
  wire[14:0] ln_if_142_acc_nl;
  wire[15:0] nl_ln_if_142_acc_nl;
  wire[11:0] ln_if_143_acc_nl;
  wire[12:0] nl_ln_if_143_acc_nl;
  wire[13:0] ln_if_141_acc_nl;
  wire[14:0] nl_ln_if_141_acc_nl;
  wire[14:0] ln_if_140_acc_nl;
  wire[15:0] nl_ln_if_140_acc_nl;
  wire[14:0] ln_if_52_acc_nl;
  wire[15:0] nl_ln_if_52_acc_nl;
  wire[14:0] ln_if_53_acc_nl;
  wire[15:0] nl_ln_if_53_acc_nl;
  wire[12:0] ln_if_49_acc_nl;
  wire[13:0] nl_ln_if_49_acc_nl;
  wire[14:0] ln_if_50_acc_nl;
  wire[15:0] nl_ln_if_50_acc_nl;
  wire[8:0] ln_if_6_acc_nl;
  wire[9:0] nl_ln_if_6_acc_nl;
  wire[5:0] ln_if_7_acc_nl;
  wire[6:0] nl_ln_if_7_acc_nl;
  wire[12:0] ln_if_139_acc_nl;
  wire[13:0] nl_ln_if_139_acc_nl;
  wire[14:0] ln_if_138_acc_nl;
  wire[15:0] nl_ln_if_138_acc_nl;
  wire[13:0] ln_if_137_acc_nl;
  wire[14:0] nl_ln_if_137_acc_nl;
  wire[14:0] ln_if_136_acc_nl;
  wire[15:0] nl_ln_if_136_acc_nl;
  wire[10:0] ln_if_135_acc_nl;
  wire[11:0] nl_ln_if_135_acc_nl;
  wire[14:0] ln_if_134_acc_nl;
  wire[15:0] nl_ln_if_134_acc_nl;
  wire[13:0] ln_if_133_acc_nl;
  wire[14:0] nl_ln_if_133_acc_nl;
  wire[14:0] ln_if_132_acc_nl;
  wire[15:0] nl_ln_if_132_acc_nl;
  wire[12:0] ln_if_131_acc_nl;
  wire[13:0] nl_ln_if_131_acc_nl;
  wire[14:0] ln_if_130_acc_nl;
  wire[15:0] nl_ln_if_130_acc_nl;
  wire[13:0] ln_if_129_acc_nl;
  wire[14:0] nl_ln_if_129_acc_nl;
  wire[14:0] ln_if_128_acc_nl;
  wire[15:0] nl_ln_if_128_acc_nl;
  wire[11:0] ln_if_127_acc_nl;
  wire[12:0] nl_ln_if_127_acc_nl;
  wire[14:0] ln_if_126_acc_nl;
  wire[15:0] nl_ln_if_126_acc_nl;
  wire[13:0] ln_if_125_acc_nl;
  wire[14:0] nl_ln_if_125_acc_nl;
  wire[14:0] ln_if_124_acc_nl;
  wire[15:0] nl_ln_if_124_acc_nl;
  wire[12:0] ln_if_123_acc_nl;
  wire[13:0] nl_ln_if_123_acc_nl;
  wire[14:0] ln_if_122_acc_nl;
  wire[15:0] nl_ln_if_122_acc_nl;
  wire[13:0] ln_if_121_acc_nl;
  wire[14:0] nl_ln_if_121_acc_nl;
  wire[14:0] ln_if_120_acc_nl;
  wire[15:0] nl_ln_if_120_acc_nl;
  wire[9:0] ln_if_119_acc_nl;
  wire[10:0] nl_ln_if_119_acc_nl;
  wire[14:0] ln_if_118_acc_nl;
  wire[15:0] nl_ln_if_118_acc_nl;
  wire[13:0] ln_if_117_acc_nl;
  wire[14:0] nl_ln_if_117_acc_nl;
  wire[14:0] ln_if_116_acc_nl;
  wire[15:0] nl_ln_if_116_acc_nl;
  wire[14:0] ln_if_115_acc_nl;
  wire[15:0] nl_ln_if_115_acc_nl;
  wire[10:0] ln_if_114_acc_nl;
  wire[11:0] nl_ln_if_114_acc_nl;
  wire[14:0] ln_if_113_acc_nl;
  wire[15:0] nl_ln_if_113_acc_nl;
  wire[13:0] ln_if_112_acc_nl;
  wire[14:0] nl_ln_if_112_acc_nl;
  wire[14:0] ln_if_111_acc_nl;
  wire[15:0] nl_ln_if_111_acc_nl;
  wire[12:0] ln_if_110_acc_nl;
  wire[13:0] nl_ln_if_110_acc_nl;
  wire[14:0] ln_if_109_acc_nl;
  wire[15:0] nl_ln_if_109_acc_nl;
  wire[14:0] ln_if_108_acc_nl;
  wire[15:0] nl_ln_if_108_acc_nl;
  wire[13:0] ln_if_107_acc_nl;
  wire[14:0] nl_ln_if_107_acc_nl;
  wire[14:0] ln_if_106_acc_nl;
  wire[15:0] nl_ln_if_106_acc_nl;
  wire[12:0] ln_if_105_acc_nl;
  wire[13:0] nl_ln_if_105_acc_nl;
  wire[14:0] ln_if_104_acc_nl;
  wire[15:0] nl_ln_if_104_acc_nl;
  wire[13:0] ln_if_103_acc_nl;
  wire[14:0] nl_ln_if_103_acc_nl;
  wire[14:0] ln_if_102_acc_nl;
  wire[15:0] nl_ln_if_102_acc_nl;
  wire[14:0] ln_if_101_acc_nl;
  wire[15:0] nl_ln_if_101_acc_nl;
  wire[12:0] ln_if_100_acc_nl;
  wire[13:0] nl_ln_if_100_acc_nl;
  wire[14:0] ln_if_99_acc_nl;
  wire[15:0] nl_ln_if_99_acc_nl;
  wire[13:0] ln_if_98_acc_nl;
  wire[14:0] nl_ln_if_98_acc_nl;
  wire[14:0] ln_if_97_acc_nl;
  wire[15:0] nl_ln_if_97_acc_nl;
  wire[11:0] ln_if_96_acc_nl;
  wire[12:0] nl_ln_if_96_acc_nl;
  wire[14:0] ln_if_95_acc_nl;
  wire[15:0] nl_ln_if_95_acc_nl;
  wire[14:0] ln_if_94_acc_nl;
  wire[15:0] nl_ln_if_94_acc_nl;
  wire[13:0] ln_if_93_acc_nl;
  wire[14:0] nl_ln_if_93_acc_nl;
  wire[14:0] ln_if_92_acc_nl;
  wire[15:0] nl_ln_if_92_acc_nl;
  wire[11:0] ln_if_91_acc_nl;
  wire[12:0] nl_ln_if_91_acc_nl;
  wire[14:0] ln_if_90_acc_nl;
  wire[15:0] nl_ln_if_90_acc_nl;
  wire[13:0] ln_if_89_acc_nl;
  wire[14:0] nl_ln_if_89_acc_nl;
  wire[14:0] ln_if_88_acc_nl;
  wire[15:0] nl_ln_if_88_acc_nl;
  wire[14:0] ln_if_87_acc_nl;
  wire[15:0] nl_ln_if_87_acc_nl;
  wire[11:0] ln_if_86_acc_nl;
  wire[12:0] nl_ln_if_86_acc_nl;
  wire[14:0] ln_if_85_acc_nl;
  wire[15:0] nl_ln_if_85_acc_nl;
  wire[13:0] ln_if_84_acc_nl;
  wire[14:0] nl_ln_if_84_acc_nl;
  wire[14:0] ln_if_83_acc_nl;
  wire[15:0] nl_ln_if_83_acc_nl;
  wire[12:0] ln_if_82_acc_nl;
  wire[13:0] nl_ln_if_82_acc_nl;
  wire[14:0] ln_if_81_acc_nl;
  wire[15:0] nl_ln_if_81_acc_nl;
  wire[14:0] ln_if_80_acc_nl;
  wire[15:0] nl_ln_if_80_acc_nl;
  wire[13:0] ln_if_79_acc_nl;
  wire[14:0] nl_ln_if_79_acc_nl;
  wire[14:0] ln_if_78_acc_nl;
  wire[15:0] nl_ln_if_78_acc_nl;
  wire[12:0] ln_if_77_acc_nl;
  wire[13:0] nl_ln_if_77_acc_nl;
  wire[14:0] ln_if_76_acc_nl;
  wire[15:0] nl_ln_if_76_acc_nl;
  wire[13:0] ln_if_75_acc_nl;
  wire[14:0] nl_ln_if_75_acc_nl;
  wire[14:0] ln_if_74_acc_nl;
  wire[15:0] nl_ln_if_74_acc_nl;
  wire[14:0] ln_if_73_acc_nl;
  wire[15:0] nl_ln_if_73_acc_nl;
  wire[12:0] ln_if_72_acc_nl;
  wire[13:0] nl_ln_if_72_acc_nl;
  wire[14:0] ln_if_71_acc_nl;
  wire[15:0] nl_ln_if_71_acc_nl;
  wire[13:0] ln_if_70_acc_nl;
  wire[14:0] nl_ln_if_70_acc_nl;
  wire[14:0] ln_if_69_acc_nl;
  wire[15:0] nl_ln_if_69_acc_nl;
  wire[8:0] ln_if_68_acc_nl;
  wire[9:0] nl_ln_if_68_acc_nl;
  wire[14:0] ln_if_67_acc_nl;
  wire[15:0] nl_ln_if_67_acc_nl;
  wire[14:0] ln_if_66_acc_nl;
  wire[15:0] nl_ln_if_66_acc_nl;
  wire[13:0] ln_if_65_acc_nl;
  wire[14:0] nl_ln_if_65_acc_nl;
  wire[14:0] ln_if_64_acc_nl;
  wire[15:0] nl_ln_if_64_acc_nl;
  wire[10:0] ln_if_63_acc_nl;
  wire[11:0] nl_ln_if_63_acc_nl;
  wire[14:0] ln_if_62_acc_nl;
  wire[15:0] nl_ln_if_62_acc_nl;
  wire[13:0] ln_if_61_acc_nl;
  wire[14:0] nl_ln_if_61_acc_nl;
  wire[14:0] ln_if_60_acc_nl;
  wire[15:0] nl_ln_if_60_acc_nl;
  wire[14:0] ln_if_59_acc_nl;
  wire[15:0] nl_ln_if_59_acc_nl;
  wire[9:0] ln_if_58_acc_nl;
  wire[10:0] nl_ln_if_58_acc_nl;
  wire[14:0] ln_if_57_acc_nl;
  wire[15:0] nl_ln_if_57_acc_nl;
  wire[13:0] ln_if_56_acc_nl;
  wire[14:0] nl_ln_if_56_acc_nl;
  wire[14:0] ln_if_55_acc_nl;
  wire[15:0] nl_ln_if_55_acc_nl;
  wire[12:0] ln_if_54_acc_nl;
  wire[13:0] nl_ln_if_54_acc_nl;
  wire[13:0] ln_if_51_acc_nl;
  wire[14:0] nl_ln_if_51_acc_nl;
  wire[14:0] ln_if_48_acc_nl;
  wire[15:0] nl_ln_if_48_acc_nl;
  wire[13:0] ln_if_47_acc_nl;
  wire[14:0] nl_ln_if_47_acc_nl;
  wire[14:0] ln_if_46_acc_nl;
  wire[15:0] nl_ln_if_46_acc_nl;
  wire[14:0] ln_if_45_acc_nl;
  wire[15:0] nl_ln_if_45_acc_nl;
  wire[12:0] ln_if_44_acc_nl;
  wire[13:0] nl_ln_if_44_acc_nl;
  wire[14:0] ln_if_43_acc_nl;
  wire[15:0] nl_ln_if_43_acc_nl;
  wire[13:0] ln_if_42_acc_nl;
  wire[14:0] nl_ln_if_42_acc_nl;
  wire[14:0] ln_if_41_acc_nl;
  wire[15:0] nl_ln_if_41_acc_nl;
  wire[11:0] ln_if_40_acc_nl;
  wire[12:0] nl_ln_if_40_acc_nl;
  wire[14:0] ln_if_39_acc_nl;
  wire[15:0] nl_ln_if_39_acc_nl;
  wire[14:0] ln_if_38_acc_nl;
  wire[15:0] nl_ln_if_38_acc_nl;
  wire[13:0] ln_if_37_acc_nl;
  wire[14:0] nl_ln_if_37_acc_nl;
  wire[14:0] ln_if_36_acc_nl;
  wire[15:0] nl_ln_if_36_acc_nl;
  wire[11:0] ln_if_35_acc_nl;
  wire[12:0] nl_ln_if_35_acc_nl;
  wire[14:0] ln_if_34_acc_nl;
  wire[15:0] nl_ln_if_34_acc_nl;
  wire[13:0] ln_if_33_acc_nl;
  wire[14:0] nl_ln_if_33_acc_nl;
  wire[14:0] ln_if_32_acc_nl;
  wire[15:0] nl_ln_if_32_acc_nl;
  wire[14:0] ln_if_31_acc_nl;
  wire[15:0] nl_ln_if_31_acc_nl;
  wire[11:0] ln_if_30_acc_nl;
  wire[12:0] nl_ln_if_30_acc_nl;
  wire[14:0] ln_if_29_acc_nl;
  wire[15:0] nl_ln_if_29_acc_nl;
  wire[13:0] ln_if_28_acc_nl;
  wire[14:0] nl_ln_if_28_acc_nl;
  wire[14:0] ln_if_27_acc_nl;
  wire[15:0] nl_ln_if_27_acc_nl;
  wire[12:0] ln_if_26_acc_nl;
  wire[13:0] nl_ln_if_26_acc_nl;
  wire[14:0] ln_if_25_acc_nl;
  wire[15:0] nl_ln_if_25_acc_nl;
  wire[14:0] ln_if_24_acc_nl;
  wire[15:0] nl_ln_if_24_acc_nl;
  wire[13:0] ln_if_23_acc_nl;
  wire[14:0] nl_ln_if_23_acc_nl;
  wire[14:0] ln_if_22_acc_nl;
  wire[15:0] nl_ln_if_22_acc_nl;
  wire[12:0] ln_if_21_acc_nl;
  wire[13:0] nl_ln_if_21_acc_nl;
  wire[14:0] ln_if_20_acc_nl;
  wire[15:0] nl_ln_if_20_acc_nl;
  wire[13:0] ln_if_19_acc_nl;
  wire[14:0] nl_ln_if_19_acc_nl;
  wire[14:0] ln_if_18_acc_nl;
  wire[15:0] nl_ln_if_18_acc_nl;
  wire[14:0] ln_if_17_acc_nl;
  wire[15:0] nl_ln_if_17_acc_nl;
  wire[12:0] ln_if_16_acc_nl;
  wire[13:0] nl_ln_if_16_acc_nl;
  wire[14:0] ln_if_15_acc_nl;
  wire[15:0] nl_ln_if_15_acc_nl;
  wire[13:0] ln_if_14_acc_nl;
  wire[14:0] nl_ln_if_14_acc_nl;
  wire[14:0] ln_if_13_acc_nl;
  wire[15:0] nl_ln_if_13_acc_nl;
  wire[10:0] ln_if_12_acc_nl;
  wire[11:0] nl_ln_if_12_acc_nl;
  wire[14:0] ln_if_11_acc_nl;
  wire[15:0] nl_ln_if_11_acc_nl;
  wire[14:0] ln_if_10_acc_nl;
  wire[15:0] nl_ln_if_10_acc_nl;
  wire[13:0] ln_if_9_acc_nl;
  wire[14:0] nl_ln_if_9_acc_nl;
  wire[14:0] ln_if_8_acc_nl;
  wire[15:0] nl_ln_if_8_acc_nl;
  wire[8:0] ln_if_4_acc_nl;
  wire[9:0] nl_ln_if_4_acc_nl;
  wire[7:0] ln_if_5_acc_nl;
  wire[8:0] nl_ln_if_5_acc_nl;
  wire[6:0] ln_if_3_acc_nl;
  wire[7:0] nl_ln_if_3_acc_nl;
  wire[8:0] ln_if_2_acc_nl;
  wire[9:0] nl_ln_if_2_acc_nl;
  wire[12:0] ln_1_if_252_acc_nl;
  wire[13:0] nl_ln_1_if_252_acc_nl;
  wire[14:0] ln_1_if_244_acc_nl;
  wire[15:0] nl_ln_1_if_244_acc_nl;
  wire[13:0] ln_1_if_245_acc_nl;
  wire[14:0] nl_ln_1_if_245_acc_nl;
  wire[10:0] ln_1_if_251_acc_nl;
  wire[11:0] nl_ln_1_if_251_acc_nl;
  wire[12:0] ln_1_if_250_acc_nl;
  wire[13:0] nl_ln_1_if_250_acc_nl;
  wire[11:0] ln_1_if_249_acc_nl;
  wire[12:0] nl_ln_1_if_249_acc_nl;
  wire[12:0] ln_1_if_248_acc_nl;
  wire[13:0] nl_ln_1_if_248_acc_nl;
  wire[9:0] ln_1_if_247_acc_nl;
  wire[10:0] nl_ln_1_if_247_acc_nl;
  wire[14:0] ln_1_if_246_acc_nl;
  wire[15:0] nl_ln_1_if_246_acc_nl;
  wire[7:0] ln_1_if_1_acc_nl;
  wire[8:0] nl_ln_1_if_1_acc_nl;
  wire[14:0] ln_1_if_144_acc_nl;
  wire[15:0] nl_ln_1_if_144_acc_nl;
  wire[13:0] ln_1_if_145_acc_nl;
  wire[14:0] nl_ln_1_if_145_acc_nl;
  wire[12:0] ln_1_if_243_acc_nl;
  wire[13:0] nl_ln_1_if_243_acc_nl;
  wire[14:0] ln_1_if_242_acc_nl;
  wire[15:0] nl_ln_1_if_242_acc_nl;
  wire[13:0] ln_1_if_241_acc_nl;
  wire[14:0] nl_ln_1_if_241_acc_nl;
  wire[14:0] ln_1_if_240_acc_nl;
  wire[15:0] nl_ln_1_if_240_acc_nl;
  wire[11:0] ln_1_if_239_acc_nl;
  wire[12:0] nl_ln_1_if_239_acc_nl;
  wire[14:0] ln_1_if_238_acc_nl;
  wire[15:0] nl_ln_1_if_238_acc_nl;
  wire[13:0] ln_1_if_237_acc_nl;
  wire[14:0] nl_ln_1_if_237_acc_nl;
  wire[14:0] ln_1_if_236_acc_nl;
  wire[15:0] nl_ln_1_if_236_acc_nl;
  wire[12:0] ln_1_if_235_acc_nl;
  wire[13:0] nl_ln_1_if_235_acc_nl;
  wire[14:0] ln_1_if_234_acc_nl;
  wire[15:0] nl_ln_1_if_234_acc_nl;
  wire[13:0] ln_1_if_233_acc_nl;
  wire[14:0] nl_ln_1_if_233_acc_nl;
  wire[14:0] ln_1_if_232_acc_nl;
  wire[15:0] nl_ln_1_if_232_acc_nl;
  wire[10:0] ln_1_if_231_acc_nl;
  wire[11:0] nl_ln_1_if_231_acc_nl;
  wire[14:0] ln_1_if_230_acc_nl;
  wire[15:0] nl_ln_1_if_230_acc_nl;
  wire[13:0] ln_1_if_229_acc_nl;
  wire[14:0] nl_ln_1_if_229_acc_nl;
  wire[14:0] ln_1_if_228_acc_nl;
  wire[15:0] nl_ln_1_if_228_acc_nl;
  wire[12:0] ln_1_if_227_acc_nl;
  wire[13:0] nl_ln_1_if_227_acc_nl;
  wire[14:0] ln_1_if_226_acc_nl;
  wire[15:0] nl_ln_1_if_226_acc_nl;
  wire[13:0] ln_1_if_225_acc_nl;
  wire[14:0] nl_ln_1_if_225_acc_nl;
  wire[14:0] ln_1_if_224_acc_nl;
  wire[15:0] nl_ln_1_if_224_acc_nl;
  wire[11:0] ln_1_if_223_acc_nl;
  wire[12:0] nl_ln_1_if_223_acc_nl;
  wire[14:0] ln_1_if_222_acc_nl;
  wire[15:0] nl_ln_1_if_222_acc_nl;
  wire[13:0] ln_1_if_221_acc_nl;
  wire[14:0] nl_ln_1_if_221_acc_nl;
  wire[14:0] ln_1_if_220_acc_nl;
  wire[15:0] nl_ln_1_if_220_acc_nl;
  wire[12:0] ln_1_if_219_acc_nl;
  wire[13:0] nl_ln_1_if_219_acc_nl;
  wire[14:0] ln_1_if_218_acc_nl;
  wire[15:0] nl_ln_1_if_218_acc_nl;
  wire[13:0] ln_1_if_217_acc_nl;
  wire[14:0] nl_ln_1_if_217_acc_nl;
  wire[14:0] ln_1_if_216_acc_nl;
  wire[15:0] nl_ln_1_if_216_acc_nl;
  wire[8:0] ln_1_if_215_acc_nl;
  wire[9:0] nl_ln_1_if_215_acc_nl;
  wire[14:0] ln_1_if_214_acc_nl;
  wire[15:0] nl_ln_1_if_214_acc_nl;
  wire[13:0] ln_1_if_213_acc_nl;
  wire[14:0] nl_ln_1_if_213_acc_nl;
  wire[14:0] ln_1_if_212_acc_nl;
  wire[15:0] nl_ln_1_if_212_acc_nl;
  wire[12:0] ln_1_if_211_acc_nl;
  wire[13:0] nl_ln_1_if_211_acc_nl;
  wire[14:0] ln_1_if_210_acc_nl;
  wire[15:0] nl_ln_1_if_210_acc_nl;
  wire[13:0] ln_1_if_209_acc_nl;
  wire[14:0] nl_ln_1_if_209_acc_nl;
  wire[14:0] ln_1_if_208_acc_nl;
  wire[15:0] nl_ln_1_if_208_acc_nl;
  wire[11:0] ln_1_if_207_acc_nl;
  wire[12:0] nl_ln_1_if_207_acc_nl;
  wire[14:0] ln_1_if_206_acc_nl;
  wire[15:0] nl_ln_1_if_206_acc_nl;
  wire[13:0] ln_1_if_205_acc_nl;
  wire[14:0] nl_ln_1_if_205_acc_nl;
  wire[14:0] ln_1_if_204_acc_nl;
  wire[15:0] nl_ln_1_if_204_acc_nl;
  wire[12:0] ln_1_if_203_acc_nl;
  wire[13:0] nl_ln_1_if_203_acc_nl;
  wire[14:0] ln_1_if_202_acc_nl;
  wire[15:0] nl_ln_1_if_202_acc_nl;
  wire[13:0] ln_1_if_201_acc_nl;
  wire[14:0] nl_ln_1_if_201_acc_nl;
  wire[14:0] ln_1_if_200_acc_nl;
  wire[15:0] nl_ln_1_if_200_acc_nl;
  wire[10:0] ln_1_if_199_acc_nl;
  wire[11:0] nl_ln_1_if_199_acc_nl;
  wire[14:0] ln_1_if_198_acc_nl;
  wire[15:0] nl_ln_1_if_198_acc_nl;
  wire[13:0] ln_1_if_197_acc_nl;
  wire[14:0] nl_ln_1_if_197_acc_nl;
  wire[14:0] ln_1_if_196_acc_nl;
  wire[15:0] nl_ln_1_if_196_acc_nl;
  wire[12:0] ln_1_if_195_acc_nl;
  wire[13:0] nl_ln_1_if_195_acc_nl;
  wire[14:0] ln_1_if_194_acc_nl;
  wire[15:0] nl_ln_1_if_194_acc_nl;
  wire[13:0] ln_1_if_193_acc_nl;
  wire[14:0] nl_ln_1_if_193_acc_nl;
  wire[14:0] ln_1_if_192_acc_nl;
  wire[15:0] nl_ln_1_if_192_acc_nl;
  wire[11:0] ln_1_if_191_acc_nl;
  wire[12:0] nl_ln_1_if_191_acc_nl;
  wire[14:0] ln_1_if_190_acc_nl;
  wire[15:0] nl_ln_1_if_190_acc_nl;
  wire[13:0] ln_1_if_189_acc_nl;
  wire[14:0] nl_ln_1_if_189_acc_nl;
  wire[14:0] ln_1_if_188_acc_nl;
  wire[15:0] nl_ln_1_if_188_acc_nl;
  wire[12:0] ln_1_if_187_acc_nl;
  wire[13:0] nl_ln_1_if_187_acc_nl;
  wire[14:0] ln_1_if_186_acc_nl;
  wire[15:0] nl_ln_1_if_186_acc_nl;
  wire[13:0] ln_1_if_185_acc_nl;
  wire[14:0] nl_ln_1_if_185_acc_nl;
  wire[14:0] ln_1_if_184_acc_nl;
  wire[15:0] nl_ln_1_if_184_acc_nl;
  wire[9:0] ln_1_if_183_acc_nl;
  wire[10:0] nl_ln_1_if_183_acc_nl;
  wire[14:0] ln_1_if_182_acc_nl;
  wire[15:0] nl_ln_1_if_182_acc_nl;
  wire[13:0] ln_1_if_181_acc_nl;
  wire[14:0] nl_ln_1_if_181_acc_nl;
  wire[14:0] ln_1_if_180_acc_nl;
  wire[15:0] nl_ln_1_if_180_acc_nl;
  wire[12:0] ln_1_if_179_acc_nl;
  wire[13:0] nl_ln_1_if_179_acc_nl;
  wire[14:0] ln_1_if_178_acc_nl;
  wire[15:0] nl_ln_1_if_178_acc_nl;
  wire[13:0] ln_1_if_177_acc_nl;
  wire[14:0] nl_ln_1_if_177_acc_nl;
  wire[14:0] ln_1_if_176_acc_nl;
  wire[15:0] nl_ln_1_if_176_acc_nl;
  wire[11:0] ln_1_if_175_acc_nl;
  wire[12:0] nl_ln_1_if_175_acc_nl;
  wire[14:0] ln_1_if_174_acc_nl;
  wire[15:0] nl_ln_1_if_174_acc_nl;
  wire[13:0] ln_1_if_173_acc_nl;
  wire[14:0] nl_ln_1_if_173_acc_nl;
  wire[14:0] ln_1_if_172_acc_nl;
  wire[15:0] nl_ln_1_if_172_acc_nl;
  wire[12:0] ln_1_if_171_acc_nl;
  wire[13:0] nl_ln_1_if_171_acc_nl;
  wire[14:0] ln_1_if_170_acc_nl;
  wire[15:0] nl_ln_1_if_170_acc_nl;
  wire[13:0] ln_1_if_169_acc_nl;
  wire[14:0] nl_ln_1_if_169_acc_nl;
  wire[14:0] ln_1_if_168_acc_nl;
  wire[15:0] nl_ln_1_if_168_acc_nl;
  wire[10:0] ln_1_if_167_acc_nl;
  wire[11:0] nl_ln_1_if_167_acc_nl;
  wire[14:0] ln_1_if_166_acc_nl;
  wire[15:0] nl_ln_1_if_166_acc_nl;
  wire[13:0] ln_1_if_165_acc_nl;
  wire[14:0] nl_ln_1_if_165_acc_nl;
  wire[14:0] ln_1_if_164_acc_nl;
  wire[15:0] nl_ln_1_if_164_acc_nl;
  wire[12:0] ln_1_if_163_acc_nl;
  wire[13:0] nl_ln_1_if_163_acc_nl;
  wire[14:0] ln_1_if_162_acc_nl;
  wire[15:0] nl_ln_1_if_162_acc_nl;
  wire[13:0] ln_1_if_161_acc_nl;
  wire[14:0] nl_ln_1_if_161_acc_nl;
  wire[14:0] ln_1_if_160_acc_nl;
  wire[15:0] nl_ln_1_if_160_acc_nl;
  wire[11:0] ln_1_if_159_acc_nl;
  wire[12:0] nl_ln_1_if_159_acc_nl;
  wire[14:0] ln_1_if_158_acc_nl;
  wire[15:0] nl_ln_1_if_158_acc_nl;
  wire[13:0] ln_1_if_157_acc_nl;
  wire[14:0] nl_ln_1_if_157_acc_nl;
  wire[14:0] ln_1_if_156_acc_nl;
  wire[15:0] nl_ln_1_if_156_acc_nl;
  wire[12:0] ln_1_if_155_acc_nl;
  wire[13:0] nl_ln_1_if_155_acc_nl;
  wire[14:0] ln_1_if_154_acc_nl;
  wire[15:0] nl_ln_1_if_154_acc_nl;
  wire[13:0] ln_1_if_153_acc_nl;
  wire[14:0] nl_ln_1_if_153_acc_nl;
  wire[14:0] ln_1_if_152_acc_nl;
  wire[15:0] nl_ln_1_if_152_acc_nl;
  wire[7:0] ln_1_if_151_acc_nl;
  wire[8:0] nl_ln_1_if_151_acc_nl;
  wire[14:0] ln_1_if_150_acc_nl;
  wire[15:0] nl_ln_1_if_150_acc_nl;
  wire[13:0] ln_1_if_149_acc_nl;
  wire[14:0] nl_ln_1_if_149_acc_nl;
  wire[14:0] ln_1_if_148_acc_nl;
  wire[15:0] nl_ln_1_if_148_acc_nl;
  wire[12:0] ln_1_if_147_acc_nl;
  wire[13:0] nl_ln_1_if_147_acc_nl;
  wire[14:0] ln_1_if_146_acc_nl;
  wire[15:0] nl_ln_1_if_146_acc_nl;
  wire[14:0] ln_1_if_142_acc_nl;
  wire[15:0] nl_ln_1_if_142_acc_nl;
  wire[11:0] ln_1_if_143_acc_nl;
  wire[12:0] nl_ln_1_if_143_acc_nl;
  wire[13:0] ln_1_if_141_acc_nl;
  wire[14:0] nl_ln_1_if_141_acc_nl;
  wire[14:0] ln_1_if_140_acc_nl;
  wire[15:0] nl_ln_1_if_140_acc_nl;
  wire[14:0] ln_1_if_52_acc_nl;
  wire[15:0] nl_ln_1_if_52_acc_nl;
  wire[14:0] ln_1_if_53_acc_nl;
  wire[15:0] nl_ln_1_if_53_acc_nl;
  wire[12:0] ln_1_if_49_acc_nl;
  wire[13:0] nl_ln_1_if_49_acc_nl;
  wire[14:0] ln_1_if_50_acc_nl;
  wire[15:0] nl_ln_1_if_50_acc_nl;
  wire[8:0] ln_1_if_6_acc_nl;
  wire[9:0] nl_ln_1_if_6_acc_nl;
  wire[5:0] ln_1_if_7_acc_nl;
  wire[6:0] nl_ln_1_if_7_acc_nl;
  wire[12:0] ln_1_if_139_acc_nl;
  wire[13:0] nl_ln_1_if_139_acc_nl;
  wire[14:0] ln_1_if_138_acc_nl;
  wire[15:0] nl_ln_1_if_138_acc_nl;
  wire[13:0] ln_1_if_137_acc_nl;
  wire[14:0] nl_ln_1_if_137_acc_nl;
  wire[14:0] ln_1_if_136_acc_nl;
  wire[15:0] nl_ln_1_if_136_acc_nl;
  wire[10:0] ln_1_if_135_acc_nl;
  wire[11:0] nl_ln_1_if_135_acc_nl;
  wire[14:0] ln_1_if_134_acc_nl;
  wire[15:0] nl_ln_1_if_134_acc_nl;
  wire[13:0] ln_1_if_133_acc_nl;
  wire[14:0] nl_ln_1_if_133_acc_nl;
  wire[14:0] ln_1_if_132_acc_nl;
  wire[15:0] nl_ln_1_if_132_acc_nl;
  wire[12:0] ln_1_if_131_acc_nl;
  wire[13:0] nl_ln_1_if_131_acc_nl;
  wire[14:0] ln_1_if_130_acc_nl;
  wire[15:0] nl_ln_1_if_130_acc_nl;
  wire[13:0] ln_1_if_129_acc_nl;
  wire[14:0] nl_ln_1_if_129_acc_nl;
  wire[14:0] ln_1_if_128_acc_nl;
  wire[15:0] nl_ln_1_if_128_acc_nl;
  wire[11:0] ln_1_if_127_acc_nl;
  wire[12:0] nl_ln_1_if_127_acc_nl;
  wire[14:0] ln_1_if_126_acc_nl;
  wire[15:0] nl_ln_1_if_126_acc_nl;
  wire[13:0] ln_1_if_125_acc_nl;
  wire[14:0] nl_ln_1_if_125_acc_nl;
  wire[14:0] ln_1_if_124_acc_nl;
  wire[15:0] nl_ln_1_if_124_acc_nl;
  wire[12:0] ln_1_if_123_acc_nl;
  wire[13:0] nl_ln_1_if_123_acc_nl;
  wire[14:0] ln_1_if_122_acc_nl;
  wire[15:0] nl_ln_1_if_122_acc_nl;
  wire[13:0] ln_1_if_121_acc_nl;
  wire[14:0] nl_ln_1_if_121_acc_nl;
  wire[14:0] ln_1_if_120_acc_nl;
  wire[15:0] nl_ln_1_if_120_acc_nl;
  wire[9:0] ln_1_if_119_acc_nl;
  wire[10:0] nl_ln_1_if_119_acc_nl;
  wire[14:0] ln_1_if_118_acc_nl;
  wire[15:0] nl_ln_1_if_118_acc_nl;
  wire[13:0] ln_1_if_117_acc_nl;
  wire[14:0] nl_ln_1_if_117_acc_nl;
  wire[14:0] ln_1_if_116_acc_nl;
  wire[15:0] nl_ln_1_if_116_acc_nl;
  wire[14:0] ln_1_if_115_acc_nl;
  wire[15:0] nl_ln_1_if_115_acc_nl;
  wire[10:0] ln_1_if_114_acc_nl;
  wire[11:0] nl_ln_1_if_114_acc_nl;
  wire[14:0] ln_1_if_113_acc_nl;
  wire[15:0] nl_ln_1_if_113_acc_nl;
  wire[13:0] ln_1_if_112_acc_nl;
  wire[14:0] nl_ln_1_if_112_acc_nl;
  wire[14:0] ln_1_if_111_acc_nl;
  wire[15:0] nl_ln_1_if_111_acc_nl;
  wire[12:0] ln_1_if_110_acc_nl;
  wire[13:0] nl_ln_1_if_110_acc_nl;
  wire[14:0] ln_1_if_109_acc_nl;
  wire[15:0] nl_ln_1_if_109_acc_nl;
  wire[14:0] ln_1_if_108_acc_nl;
  wire[15:0] nl_ln_1_if_108_acc_nl;
  wire[13:0] ln_1_if_107_acc_nl;
  wire[14:0] nl_ln_1_if_107_acc_nl;
  wire[14:0] ln_1_if_106_acc_nl;
  wire[15:0] nl_ln_1_if_106_acc_nl;
  wire[12:0] ln_1_if_105_acc_nl;
  wire[13:0] nl_ln_1_if_105_acc_nl;
  wire[14:0] ln_1_if_104_acc_nl;
  wire[15:0] nl_ln_1_if_104_acc_nl;
  wire[13:0] ln_1_if_103_acc_nl;
  wire[14:0] nl_ln_1_if_103_acc_nl;
  wire[14:0] ln_1_if_102_acc_nl;
  wire[15:0] nl_ln_1_if_102_acc_nl;
  wire[14:0] ln_1_if_101_acc_nl;
  wire[15:0] nl_ln_1_if_101_acc_nl;
  wire[12:0] ln_1_if_100_acc_nl;
  wire[13:0] nl_ln_1_if_100_acc_nl;
  wire[14:0] ln_1_if_99_acc_nl;
  wire[15:0] nl_ln_1_if_99_acc_nl;
  wire[13:0] ln_1_if_98_acc_nl;
  wire[14:0] nl_ln_1_if_98_acc_nl;
  wire[14:0] ln_1_if_97_acc_nl;
  wire[15:0] nl_ln_1_if_97_acc_nl;
  wire[11:0] ln_1_if_96_acc_nl;
  wire[12:0] nl_ln_1_if_96_acc_nl;
  wire[14:0] ln_1_if_95_acc_nl;
  wire[15:0] nl_ln_1_if_95_acc_nl;
  wire[14:0] ln_1_if_94_acc_nl;
  wire[15:0] nl_ln_1_if_94_acc_nl;
  wire[13:0] ln_1_if_93_acc_nl;
  wire[14:0] nl_ln_1_if_93_acc_nl;
  wire[14:0] ln_1_if_92_acc_nl;
  wire[15:0] nl_ln_1_if_92_acc_nl;
  wire[11:0] ln_1_if_91_acc_nl;
  wire[12:0] nl_ln_1_if_91_acc_nl;
  wire[14:0] ln_1_if_90_acc_nl;
  wire[15:0] nl_ln_1_if_90_acc_nl;
  wire[13:0] ln_1_if_89_acc_nl;
  wire[14:0] nl_ln_1_if_89_acc_nl;
  wire[14:0] ln_1_if_88_acc_nl;
  wire[15:0] nl_ln_1_if_88_acc_nl;
  wire[14:0] ln_1_if_87_acc_nl;
  wire[15:0] nl_ln_1_if_87_acc_nl;
  wire[11:0] ln_1_if_86_acc_nl;
  wire[12:0] nl_ln_1_if_86_acc_nl;
  wire[14:0] ln_1_if_85_acc_nl;
  wire[15:0] nl_ln_1_if_85_acc_nl;
  wire[13:0] ln_1_if_84_acc_nl;
  wire[14:0] nl_ln_1_if_84_acc_nl;
  wire[14:0] ln_1_if_83_acc_nl;
  wire[15:0] nl_ln_1_if_83_acc_nl;
  wire[12:0] ln_1_if_82_acc_nl;
  wire[13:0] nl_ln_1_if_82_acc_nl;
  wire[14:0] ln_1_if_81_acc_nl;
  wire[15:0] nl_ln_1_if_81_acc_nl;
  wire[14:0] ln_1_if_80_acc_nl;
  wire[15:0] nl_ln_1_if_80_acc_nl;
  wire[13:0] ln_1_if_79_acc_nl;
  wire[14:0] nl_ln_1_if_79_acc_nl;
  wire[14:0] ln_1_if_78_acc_nl;
  wire[15:0] nl_ln_1_if_78_acc_nl;
  wire[12:0] ln_1_if_77_acc_nl;
  wire[13:0] nl_ln_1_if_77_acc_nl;
  wire[14:0] ln_1_if_76_acc_nl;
  wire[15:0] nl_ln_1_if_76_acc_nl;
  wire[13:0] ln_1_if_75_acc_nl;
  wire[14:0] nl_ln_1_if_75_acc_nl;
  wire[14:0] ln_1_if_74_acc_nl;
  wire[15:0] nl_ln_1_if_74_acc_nl;
  wire[14:0] ln_1_if_73_acc_nl;
  wire[15:0] nl_ln_1_if_73_acc_nl;
  wire[12:0] ln_1_if_72_acc_nl;
  wire[13:0] nl_ln_1_if_72_acc_nl;
  wire[14:0] ln_1_if_71_acc_nl;
  wire[15:0] nl_ln_1_if_71_acc_nl;
  wire[13:0] ln_1_if_70_acc_nl;
  wire[14:0] nl_ln_1_if_70_acc_nl;
  wire[14:0] ln_1_if_69_acc_nl;
  wire[15:0] nl_ln_1_if_69_acc_nl;
  wire[8:0] ln_1_if_68_acc_nl;
  wire[9:0] nl_ln_1_if_68_acc_nl;
  wire[14:0] ln_1_if_67_acc_nl;
  wire[15:0] nl_ln_1_if_67_acc_nl;
  wire[14:0] ln_1_if_66_acc_nl;
  wire[15:0] nl_ln_1_if_66_acc_nl;
  wire[13:0] ln_1_if_65_acc_nl;
  wire[14:0] nl_ln_1_if_65_acc_nl;
  wire[14:0] ln_1_if_64_acc_nl;
  wire[15:0] nl_ln_1_if_64_acc_nl;
  wire[10:0] ln_1_if_63_acc_nl;
  wire[11:0] nl_ln_1_if_63_acc_nl;
  wire[14:0] ln_1_if_62_acc_nl;
  wire[15:0] nl_ln_1_if_62_acc_nl;
  wire[13:0] ln_1_if_61_acc_nl;
  wire[14:0] nl_ln_1_if_61_acc_nl;
  wire[14:0] ln_1_if_60_acc_nl;
  wire[15:0] nl_ln_1_if_60_acc_nl;
  wire[14:0] ln_1_if_59_acc_nl;
  wire[15:0] nl_ln_1_if_59_acc_nl;
  wire[9:0] ln_1_if_58_acc_nl;
  wire[10:0] nl_ln_1_if_58_acc_nl;
  wire[14:0] ln_1_if_57_acc_nl;
  wire[15:0] nl_ln_1_if_57_acc_nl;
  wire[13:0] ln_1_if_56_acc_nl;
  wire[14:0] nl_ln_1_if_56_acc_nl;
  wire[14:0] ln_1_if_55_acc_nl;
  wire[15:0] nl_ln_1_if_55_acc_nl;
  wire[12:0] ln_1_if_54_acc_nl;
  wire[13:0] nl_ln_1_if_54_acc_nl;
  wire[13:0] ln_1_if_51_acc_nl;
  wire[14:0] nl_ln_1_if_51_acc_nl;
  wire[14:0] ln_1_if_48_acc_nl;
  wire[15:0] nl_ln_1_if_48_acc_nl;
  wire[13:0] ln_1_if_47_acc_nl;
  wire[14:0] nl_ln_1_if_47_acc_nl;
  wire[14:0] ln_1_if_46_acc_nl;
  wire[15:0] nl_ln_1_if_46_acc_nl;
  wire[14:0] ln_1_if_45_acc_nl;
  wire[15:0] nl_ln_1_if_45_acc_nl;
  wire[12:0] ln_1_if_44_acc_nl;
  wire[13:0] nl_ln_1_if_44_acc_nl;
  wire[14:0] ln_1_if_43_acc_nl;
  wire[15:0] nl_ln_1_if_43_acc_nl;
  wire[13:0] ln_1_if_42_acc_nl;
  wire[14:0] nl_ln_1_if_42_acc_nl;
  wire[14:0] ln_1_if_41_acc_nl;
  wire[15:0] nl_ln_1_if_41_acc_nl;
  wire[11:0] ln_1_if_40_acc_nl;
  wire[12:0] nl_ln_1_if_40_acc_nl;
  wire[14:0] ln_1_if_39_acc_nl;
  wire[15:0] nl_ln_1_if_39_acc_nl;
  wire[14:0] ln_1_if_38_acc_nl;
  wire[15:0] nl_ln_1_if_38_acc_nl;
  wire[13:0] ln_1_if_37_acc_nl;
  wire[14:0] nl_ln_1_if_37_acc_nl;
  wire[14:0] ln_1_if_36_acc_nl;
  wire[15:0] nl_ln_1_if_36_acc_nl;
  wire[11:0] ln_1_if_35_acc_nl;
  wire[12:0] nl_ln_1_if_35_acc_nl;
  wire[14:0] ln_1_if_34_acc_nl;
  wire[15:0] nl_ln_1_if_34_acc_nl;
  wire[13:0] ln_1_if_33_acc_nl;
  wire[14:0] nl_ln_1_if_33_acc_nl;
  wire[14:0] ln_1_if_32_acc_nl;
  wire[15:0] nl_ln_1_if_32_acc_nl;
  wire[14:0] ln_1_if_31_acc_nl;
  wire[15:0] nl_ln_1_if_31_acc_nl;
  wire[11:0] ln_1_if_30_acc_nl;
  wire[12:0] nl_ln_1_if_30_acc_nl;
  wire[14:0] ln_1_if_29_acc_nl;
  wire[15:0] nl_ln_1_if_29_acc_nl;
  wire[13:0] ln_1_if_28_acc_nl;
  wire[14:0] nl_ln_1_if_28_acc_nl;
  wire[14:0] ln_1_if_27_acc_nl;
  wire[15:0] nl_ln_1_if_27_acc_nl;
  wire[12:0] ln_1_if_26_acc_nl;
  wire[13:0] nl_ln_1_if_26_acc_nl;
  wire[14:0] ln_1_if_25_acc_nl;
  wire[15:0] nl_ln_1_if_25_acc_nl;
  wire[14:0] ln_1_if_24_acc_nl;
  wire[15:0] nl_ln_1_if_24_acc_nl;
  wire[13:0] ln_1_if_23_acc_nl;
  wire[14:0] nl_ln_1_if_23_acc_nl;
  wire[14:0] ln_1_if_22_acc_nl;
  wire[15:0] nl_ln_1_if_22_acc_nl;
  wire[12:0] ln_1_if_21_acc_nl;
  wire[13:0] nl_ln_1_if_21_acc_nl;
  wire[14:0] ln_1_if_20_acc_nl;
  wire[15:0] nl_ln_1_if_20_acc_nl;
  wire[13:0] ln_1_if_19_acc_nl;
  wire[14:0] nl_ln_1_if_19_acc_nl;
  wire[14:0] ln_1_if_18_acc_nl;
  wire[15:0] nl_ln_1_if_18_acc_nl;
  wire[14:0] ln_1_if_17_acc_nl;
  wire[15:0] nl_ln_1_if_17_acc_nl;
  wire[12:0] ln_1_if_16_acc_nl;
  wire[13:0] nl_ln_1_if_16_acc_nl;
  wire[14:0] ln_1_if_15_acc_nl;
  wire[15:0] nl_ln_1_if_15_acc_nl;
  wire[13:0] ln_1_if_14_acc_nl;
  wire[14:0] nl_ln_1_if_14_acc_nl;
  wire[14:0] ln_1_if_13_acc_nl;
  wire[15:0] nl_ln_1_if_13_acc_nl;
  wire[10:0] ln_1_if_12_acc_nl;
  wire[11:0] nl_ln_1_if_12_acc_nl;
  wire[14:0] ln_1_if_11_acc_nl;
  wire[15:0] nl_ln_1_if_11_acc_nl;
  wire[14:0] ln_1_if_10_acc_nl;
  wire[15:0] nl_ln_1_if_10_acc_nl;
  wire[13:0] ln_1_if_9_acc_nl;
  wire[14:0] nl_ln_1_if_9_acc_nl;
  wire[14:0] ln_1_if_8_acc_nl;
  wire[15:0] nl_ln_1_if_8_acc_nl;
  wire[8:0] ln_1_if_4_acc_nl;
  wire[9:0] nl_ln_1_if_4_acc_nl;
  wire[7:0] ln_1_if_5_acc_nl;
  wire[8:0] nl_ln_1_if_5_acc_nl;
  wire[6:0] ln_1_if_3_acc_nl;
  wire[7:0] nl_ln_1_if_3_acc_nl;
  wire[8:0] ln_1_if_2_acc_nl;
  wire[9:0] nl_ln_1_if_2_acc_nl;
  wire mux_1315_nl;
  wire mux_1320_nl;
  wire mux_1326_nl;
  wire mux_1335_nl;
  wire mux_1356_nl;
  wire mux_1361_nl;
  wire or_209_nl;
  wire mux_1360_nl;
  wire or_207_nl;
  wire mux_1408_nl;
  wire mux_1416_nl;
  wire mux_1415_nl;
  wire mux_1414_nl;
  wire mux_1413_nl;
  wire mux_1412_nl;
  wire mux_1411_nl;
  wire mux_1410_nl;
  wire mux_1425_nl;
  wire mux_1424_nl;
  wire mux_1423_nl;
  wire mux_1422_nl;
  wire mux_1421_nl;
  wire mux_1431_nl;
  wire or_335_nl;
  wire mux_1434_nl;
  wire mux_1433_nl;
  wire mux_1437_nl;
  wire mux_1436_nl;
  wire or_339_nl;
  wire or_342_nl;
  wire mux_1442_nl;
  wire mux_1441_nl;
  wire mux_1440_nl;
  wire nand_117_nl;
  wire mux_1448_nl;
  wire mux_1447_nl;
  wire mux_1446_nl;
  wire nand_118_nl;
  wire or_350_nl;
  wire or_349_nl;
  wire mux_1455_nl;
  wire mux_1457_nl;
  wire nand_71_nl;
  wire mux_1468_nl;
  wire mux_1467_nl;
  wire or_359_nl;
  wire nor_189_nl;
  wire mux_1474_nl;
  wire mux_1473_nl;
  wire mux_1472_nl;
  wire or_367_nl;
  wire mux_1471_nl;
  wire mux_1479_nl;
  wire mux_1478_nl;
  wire and_308_nl;
  wire or_378_nl;
  wire or_380_nl;
  wire or_382_nl;
  wire mux_1495_nl;
  wire mux_1494_nl;
  wire mux_1493_nl;
  wire mux_1492_nl;
  wire mux_1491_nl;
  wire mux_1505_nl;
  wire mux_1504_nl;
  wire mux_1503_nl;
  wire mux_1502_nl;
  wire nand_123_nl;
  wire or_393_nl;
  wire mux_1517_nl;
  wire mux_1516_nl;
  wire or_395_nl;
  wire mux_1520_nl;
  wire mux_1519_nl;
  wire mux_1515_nl;
  wire mux_1514_nl;
  wire nand_126_nl;
  wire mux_1525_nl;
  wire and_319_nl;
  wire mux_1535_nl;
  wire mux_1534_nl;
  wire mux_1533_nl;
  wire nor_192_nl;
  wire mux_1532_nl;
  wire mux_1531_nl;
  wire mux_1530_nl;
  wire mux_1529_nl;
  wire mux_1528_nl;
  wire mux_1527_nl;
  wire or_405_nl;
  wire mux_1545_nl;
  wire mux_1544_nl;
  wire or_408_nl;
  wire mux_1543_nl;
  wire mux_1549_nl;
  wire or_411_nl;
  wire or_410_nl;
  wire mux_1563_nl;
  wire mux_1562_nl;
  wire mux_1561_nl;
  wire mux_1560_nl;
  wire mux_1559_nl;
  wire and_324_nl;
  wire mux_1557_nl;
  wire mux_1556_nl;
  wire nand_129_nl;
  wire or_421_nl;
  wire mux_1576_nl;
  wire or_426_nl;
  wire mux_1575_nl;
  wire mux_1574_nl;
  wire nand_77_nl;
  wire mux_1573_nl;
  wire or_424_nl;
  wire mux_1591_nl;
  wire or_432_nl;
  wire mux_1590_nl;
  wire mux_1589_nl;
  wire mux_1588_nl;
  wire mux_1587_nl;
  wire mux_1586_nl;
  wire mux_1585_nl;
  wire mux_1584_nl;
  wire or_441_nl;
  wire mux_1603_nl;
  wire mux_1602_nl;
  wire and_255_nl;
  wire mux_1606_nl;
  wire mux_1605_nl;
  wire mux_1601_nl;
  wire mux_1600_nl;
  wire or_445_nl;
  wire or_452_nl;
  wire mux_1610_nl;
  wire or_450_nl;
  wire mux_1620_nl;
  wire mux_1619_nl;
  wire mux_1618_nl;
  wire mux_1617_nl;
  wire mux_1616_nl;
  wire or_455_nl;
  wire mux_1615_nl;
  wire mux_1614_nl;
  wire mux_1613_nl;
  wire mux_1612_nl;
  wire mux_1626_nl;
  wire mux_1629_nl;
  wire nand_137_nl;
  wire mux_1637_nl;
  wire mux_1636_nl;
  wire mux_1635_nl;
  wire mux_1634_nl;
  wire mux_1633_nl;
  wire mux_1642_nl;
  wire mux_1651_nl;
  wire mux_1650_nl;
  wire mux_1649_nl;
  wire mux_1648_nl;
  wire mux_1647_nl;
  wire mux_1646_nl;
  wire mux_1658_nl;
  wire or_476_nl;
  wire or_474_nl;
  wire mux_1657_nl;
  wire mux_1661_nl;
  wire mux_1660_nl;
  wire or_613_nl;
  wire nand_139_nl;
  wire mux_1662_nl;
  wire mux_1668_nl;
  wire mux_1667_nl;
  wire mux_1666_nl;
  wire nor_195_nl;
  wire or_488_nl;
  wire mux_1678_nl;
  wire mux_1677_nl;
  wire mux_1676_nl;
  wire mux_1690_nl;
  wire mux_1689_nl;
  wire mux_1688_nl;
  wire mux_1687_nl;
  wire mux_1686_nl;
  wire mux_1685_nl;
  wire mux_1684_nl;
  wire mux_1683_nl;
  wire mux_1696_nl;
  wire nor_196_nl;
  wire or_506_nl;
  wire mux_1699_nl;
  wire mux_1697_nl;
  wire mux_1706_nl;
  wire nand_145_nl;
  wire mux_1705_nl;
  wire or_510_nl;
  wire mux_1704_nl;
  wire mux_1702_nl;
  wire mux_1701_nl;
  wire mux_1713_nl;
  wire mux_1712_nl;
  wire mux_1711_nl;
  wire nor_197_nl;
  wire mux_1720_nl;
  wire nor_198_nl;
  wire or_519_nl;
  wire mux_1722_nl;
  wire mux_1719_nl;
  wire and_352_nl;
  wire mux_1728_nl;
  wire mux_1734_nl;
  wire mux_1733_nl;
  wire mux_1732_nl;
  wire mux_1731_nl;
  wire mux_1730_nl;
  wire mux_1737_nl;
  wire mux_1736_nl;
  wire mux_1745_nl;
  wire mux_1744_nl;
  wire mux_1743_nl;
  wire mux_1742_nl;
  wire and_359_nl;
  wire mux_1741_nl;
  wire and_360_nl;
  wire mux_1752_nl;
  wire mux_1751_nl;
  wire mux_1755_nl;
  wire mux_1754_nl;
  wire mux_1779_nl;
  wire mux_1778_nl;
  wire mux_1777_nl;
  wire mux_1776_nl;
  wire mux_1775_nl;
  wire mux_1774_nl;
  wire mux_1773_nl;
  wire nor_205_nl;
  wire nor_206_nl;
  wire nand_84_nl;
  wire mux_1836_nl;
  wire mux_1835_nl;
  wire mux_1834_nl;
  wire mux_1833_nl;
  wire mux_1832_nl;
  wire mux_1831_nl;
  wire mux_1830_nl;
  wire mux_1850_nl;
  wire mux_1849_nl;
  wire mux_1848_nl;
  wire and_262_nl;
  wire mux_1861_nl;
  wire mux_1860_nl;
  wire mux_1771_nl;
  wire mux_1770_nl;
  wire nor_187_nl;
  wire nor_188_nl;
  wire or_548_nl;
  wire[1:0] mux_1876_nl;
  wire not_1767_nl;
  wire[11:0] if_4_for_and_19_nl;
  wire if_4_for_if_4_for_nand_6_nl;

  // Interconnect Declarations for Component Instantiations 
  ccs_out_v1 #(.rscid(32'sd1),
  .width(32'sd1)) is_random_rsci (
      .idat(is_random_rsci_idat),
      .dat(is_random_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd2),
  .width(32'sd1)) valid_rsci (
      .idat(valid_rsci_idat),
      .dat(valid_rsc_dat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd1)) epsilon_rsci (
      .dat(epsilon_rsc_dat),
      .idat(epsilon_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) is_random_triosy_obj (
      .ld(reg_is_random_triosy_obj_ld_cse),
      .lz(is_random_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) valid_triosy_obj (
      .ld(reg_is_random_triosy_obj_ld_cse),
      .lz(valid_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) epsilon_triosy_obj (
      .ld(epsilon_triosy_obj_ld),
      .lz(epsilon_triosy_lz)
    );
  assign and_276_cse = (count_sva==10'b1111111111);
  assign or_325_cse = (skip_sva_1_1_0_1!=2'b00);
  assign or_324_cse = reg_skip_ftd | (reg_skip_ftd_1!=2'b00);
  assign nand_101_cse = ~((j_lpi_1_dfm_1_3_0[3:2]==2'b11));
  assign nand_49_cse = ~((j_1_3_0_lpi_1_dfm_2_0_1[2]) & if_4_for_and_stg_1_0_sva_1);
  assign or_297_tmp = (nand_49_cse & nor_cse_1) | and_55_cse_1;
  assign nor_149_cse = ~((skip_sva_1_1_0_1[0]) | (~ first_sva));
  assign or_546_cse = shift_reg_1_sva_0 | or_tmp_306;
  assign nand_50_cse = ~((j_1_3_0_lpi_1_dfm_2_0_1[2]) & if_4_for_and_stg_1_1_sva_1);
  assign or_299_tmp = (nand_50_cse & nor_cse_1) | and_55_cse_1;
  assign or_301_tmp = (((j_1_3_0_lpi_1_dfm_2_0_1[2]) | (~ if_4_for_and_stg_1_1_sva_1))
      & nor_cse_1) | and_55_cse_1;
  assign nor_159_cse = ~((skip_sva_1_1_0_1!=2'b00) | (~ first_sva));
  assign nand_51_cse = ~((j_1_3_0_lpi_1_dfm_2_0_1[2]) & if_4_for_and_stg_1_2_sva_1);
  assign or_303_tmp = (nand_51_cse & nor_cse_1) | and_55_cse_1;
  assign or_305_tmp = (((j_1_3_0_lpi_1_dfm_2_0_1[2]) | (~ if_4_for_and_stg_1_2_sva_1))
      & nor_cse_1) | and_55_cse_1;
  assign nand_86_cse = ~(shift_reg_1_sva_0 & (~ or_tmp_356));
  assign nand_52_cse = ~((j_1_3_0_lpi_1_dfm_2_0_1[2]) & if_4_for_and_stg_1_3_sva_1);
  assign or_307_tmp = (nand_52_cse & nor_cse_1) | and_55_cse_1;
  assign and_294_cse = epsilon_rsci_idat & (count_sva==10'b1111111111);
  assign or_309_tmp = (((j_1_3_0_lpi_1_dfm_2_0_1[2]) | (~ if_4_for_and_stg_1_3_sva_1))
      & nor_cse_1) | and_55_cse_1;
  assign skip_static_init_or_ssc = (or_psp_mx0 & or_2_tmp) | and_91_tmp_1;
  assign nand_112_cse = ~((if_4_for_1_acc_tmp[4]) & (j_1_3_0_sva_2[3]));
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_38_cse = (~((~(or_dcpl_3 & (~
      (j_1_3_0_sva_2[3])))) & (if_4_for_1_acc_tmp[4]))) & (if_4_for_mux_50_tmp[9])
      & (~ nand_tmp) & (~(or_dcpl_188 | or_dcpl_185 | (if_4_for_mux_50_tmp[8:5]!=4'b1111)
      | nor_47_cse));
  assign and_298_cse = (asn_sft_lpi_1_dfm_st_1==10'b1111111111);
  assign nl_if_4_acc_1_nl = conv_s2s_15_16(if_4_acc_psp_sva_1) + 16'b1111110100111001;
  assign if_4_acc_1_nl = nl_if_4_acc_1_nl[15:0];
  assign if_4_acc_1_itm_15_1 = readslicef_16_1_15(if_4_acc_1_nl);
  assign ln_land_251_lpi_1_dfm_1_1 = ln_if_250_acc_itm_12_1 & (~ ln_if_251_acc_itm_10_1);
  assign ln_land_252_lpi_1_dfm_1_1 = ln_if_251_acc_itm_10_1 & (~ ln_if_252_acc_itm_12_1);
  assign ln_nor_9_cse_1 = ~(ln_and_248_ssc_1 | ln_if_253_acc_cse_11_sva_1);
  assign ln_nor_10_cse_1 = ~(ln_and_240_ssc_1 | ln_and_377_ssc_1 | ln_and_242_ssc_1
      | ln_and_407_ssc_1 | ln_and_244_ssc_1 | ln_and_379_ssc_1);
  assign ln_and_246_ssc_1 = ln_land_251_lpi_1_dfm_1 & (~ ln_land_252_lpi_1_dfm_1);
  assign nl_ln_if_253_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:3])
      + 12'b111111111111;
  assign ln_if_253_acc_nl = nl_ln_if_253_acc_nl[11:0];
  assign ln_if_253_acc_itm_11_1 = readslicef_12_1_11(ln_if_253_acc_nl);
  assign ln_land_248_lpi_1_dfm_1 = ln_if_247_acc_itm_9_1 & (~ ln_if_248_acc_itm_12_1);
  assign ln_land_249_lpi_1_dfm_1 = ln_if_248_acc_itm_12_1 & (~ ln_if_249_acc_itm_11_1);
  assign ln_land_250_lpi_1_dfm_1 = ln_if_249_acc_itm_11_1 & (~ ln_if_250_acc_itm_12_1);
  assign ln_and_240_ssc_1_1 = ln_if_244_acc_itm_14_1 & (~ ln_if_245_acc_itm_13_1)
      & (~(ln_land_247_lpi_1_dfm_1 | ln_land_248_lpi_1_dfm_1)) & (~(ln_land_249_lpi_1_dfm_1
      | ln_land_250_lpi_1_dfm_1)) & (~(ln_land_251_lpi_1_dfm_1_1 | ln_land_252_lpi_1_dfm_1_1));
  assign ln_land_246_lpi_1_dfm_1 = ln_if_245_acc_itm_13_1 & (~ ln_if_246_acc_itm_14_1);
  assign ln_land_247_lpi_1_dfm_1 = ln_if_246_acc_itm_14_1 & (~ ln_if_247_acc_itm_9_1);
  assign operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1 = MUX_v_14_8_2(({P1_0_1_23_10_sva_dfm_3_13_12
      , P1_0_1_23_10_sva_dfm_3_11_0}), P1_1_1_23_10_sva_dfm_3, P1_2_1_23_10_sva_dfm_3,
      P1_3_1_23_10_sva_dfm_3, P1_4_1_23_10_sva_dfm_3, P1_5_1_23_10_sva_dfm_3, P1_6_1_23_10_sva_dfm_3,
      P1_7_1_23_10_sva_dfm_3, j_1_3_0_lpi_1_dfm_2_0_1);
  assign nl_operator_24_14_false_AC_TRN_AC_WRAP_acc_nl = ({1'b1 , (~ operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)})
      + 15'b000000000000001;
  assign operator_24_14_false_AC_TRN_AC_WRAP_acc_nl = nl_operator_24_14_false_AC_TRN_AC_WRAP_acc_nl[14:0];
  assign operator_24_14_false_AC_TRN_AC_WRAP_acc_itm_14_1 = readslicef_15_1_14(operator_24_14_false_AC_TRN_AC_WRAP_acc_nl);
  assign ln_1_land_251_lpi_1_dfm_1_1 = ln_1_if_250_acc_itm_12_1 & (~ ln_1_if_251_acc_itm_10_1);
  assign ln_1_land_252_lpi_1_dfm_1_1 = ln_1_if_251_acc_itm_10_1 & (~ ln_1_if_252_acc_itm_12_1);
  assign ln_1_nor_9_cse_1 = ~(ln_1_and_248_ssc_1 | ln_1_if_253_acc_cse_11_sva_1);
  assign ln_1_nor_10_cse_1 = ~(ln_1_and_240_ssc_1 | ln_1_and_377_ssc_1 | ln_1_and_242_ssc_1
      | ln_1_and_407_ssc_1 | ln_1_and_244_ssc_1 | ln_1_and_379_ssc_1);
  assign ln_1_and_246_ssc_1 = ln_1_land_251_lpi_1_dfm_1 & (~ ln_1_land_252_lpi_1_dfm_1);
  assign nl_ln_1_if_253_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:3])
      + 12'b111111111111;
  assign ln_1_if_253_acc_nl = nl_ln_1_if_253_acc_nl[11:0];
  assign ln_1_if_253_acc_itm_11_1 = readslicef_12_1_11(ln_1_if_253_acc_nl);
  assign ln_1_land_248_lpi_1_dfm_1 = ln_1_if_247_acc_itm_9_1 & (~ ln_1_if_248_acc_itm_12_1);
  assign ln_1_land_249_lpi_1_dfm_1 = ln_1_if_248_acc_itm_12_1 & (~ ln_1_if_249_acc_itm_11_1);
  assign ln_1_land_250_lpi_1_dfm_1 = ln_1_if_249_acc_itm_11_1 & (~ ln_1_if_250_acc_itm_12_1);
  assign ln_1_and_240_ssc_1_1 = ln_1_if_244_acc_itm_14_1 & (~ ln_1_if_245_acc_itm_13_1)
      & (~(ln_1_land_247_lpi_1_dfm_1 | ln_1_land_248_lpi_1_dfm_1)) & (~(ln_1_land_249_lpi_1_dfm_1
      | ln_1_land_250_lpi_1_dfm_1)) & (~(ln_1_land_251_lpi_1_dfm_1_1 | ln_1_land_252_lpi_1_dfm_1_1));
  assign ln_1_land_246_lpi_1_dfm_1 = ln_1_if_245_acc_itm_13_1 & (~ ln_1_if_246_acc_itm_14_1);
  assign ln_1_land_247_lpi_1_dfm_1 = ln_1_if_246_acc_itm_14_1 & (~ ln_1_if_247_acc_itm_9_1);
  assign operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1
      = MUX_v_14_16_2(P2_0_1_23_10_sva_dfm_3, P2_1_1_23_10_sva_dfm_3, P2_2_1_23_10_sva_dfm_3,
      P2_3_1_23_10_sva_dfm_3, P2_4_1_23_10_sva_dfm_3, P2_5_1_23_10_sva_dfm_3, P2_6_1_23_10_sva_dfm_3,
      P2_7_1_23_10_sva_dfm_3, P2_8_1_23_10_sva_dfm_3, P2_9_1_23_10_sva_dfm_3, P2_10_1_23_10_sva_dfm_3,
      P2_11_1_23_10_sva_dfm_3, P2_12_1_23_10_sva_dfm_3, P2_13_1_23_10_sva_dfm_3,
      P2_14_1_23_10_sva_dfm_3, P2_15_1_23_10_sva_dfm_3, j_lpi_1_dfm_3_0_1);
  assign if_4_acc_psp_sva_1 = $signed((sum1_1_lpi_1_dfm_2_mx0[23:10])) - $signed((sum2_1_lpi_1_dfm_1_mx0[23:10]));
  assign ln_ln_ln_and_4_nl = (~(ln_land_251_lpi_1_dfm_1 | ln_land_252_lpi_1_dfm_1))
      & ln_nor_9_cse_1;
  assign ln_ln_ln_or_20_nl = (ln_ln_mux1h_118_psp_1_12 & ln_nor_10_cse_1) | ln_and_246_ssc_1
      | ln_land_252_lpi_1_dfm_1 | ln_and_248_ssc_1 | ln_if_253_acc_cse_11_sva_1;
  assign ln_ln_ln_or_21_nl = (~((~((ln_ln_mux1h_118_psp_1_11 & ln_nor_10_cse_1) |
      ln_and_246_ssc_1 | ln_land_252_lpi_1_dfm_1)) | ln_if_253_acc_cse_11_sva_1))
      | ln_and_248_ssc_1;
  assign ln_ln_ln_and_5_nl = ((ln_ln_mux1h_118_psp_1_10 & (~(ln_and_407_ssc_1 | ln_and_244_ssc_1
      | ln_and_379_ssc_1))) | ln_and_240_ssc_1 | ln_and_377_ssc_1 | ln_and_242_ssc_1
      | ln_and_246_ssc_1 | ln_land_252_lpi_1_dfm_1) & ln_nor_9_cse_1;
  assign ln_ln_ln_or_24_nl = (~((~(ln_and_427_itm_1 | ln_and_407_ssc_1 | ln_and_246_ssc_1))
      | ln_and_248_ssc_1)) | ln_if_253_acc_cse_11_sva_1;
  assign ln_ln_ln_or_26_nl = (ln_ln_mux1h_118_psp_1_8 & (~(ln_and_240_ssc_1 | ln_and_377_ssc_1
      | ln_and_242_ssc_1 | ln_and_379_ssc_1 | ln_and_246_ssc_1 | ln_land_252_lpi_1_dfm_1)))
      | ln_and_407_ssc_1 | ln_and_244_ssc_1 | ln_and_248_ssc_1 | ln_if_253_acc_cse_11_sva_1;
  assign ln_ln_ln_or_27_nl = (~((~((ln_ln_mux1h_118_psp_1_7 & (~(ln_and_242_ssc_1
      | ln_and_407_ssc_1 | ln_land_252_lpi_1_dfm_1))) | ln_and_240_ssc_1 | ln_and_377_ssc_1
      | ln_and_244_ssc_1 | ln_and_379_ssc_1 | ln_and_246_ssc_1)) | ln_and_248_ssc_1))
      | ln_if_253_acc_cse_11_sva_1;
  assign ln_ln_ln_and_6_nl = ((ln_ln_mux1h_118_psp_1_6 & (~(ln_and_377_ssc_1 | ln_and_407_ssc_1
      | ln_and_379_ssc_1 | ln_and_246_ssc_1))) | ln_and_240_ssc_1 | ln_and_242_ssc_1
      | ln_and_244_ssc_1 | ln_land_252_lpi_1_dfm_1) & ln_nor_9_cse_1;
  assign ln_ln_ln_or_30_nl = (ln_ln_mux1h_118_psp_1_5 & (~(ln_and_240_ssc_1 | ln_and_377_ssc_1
      | ln_and_242_ssc_1 | ln_and_379_ssc_1))) | ln_and_407_ssc_1 | ln_and_244_ssc_1
      | ln_and_246_ssc_1 | ln_land_252_lpi_1_dfm_1 | ln_and_248_ssc_1 | ln_if_253_acc_cse_11_sva_1;
  assign ln_ln_ln_and_7_nl = ((ln_ln_mux1h_118_psp_1_4 & (~(ln_and_240_ssc_1 | ln_and_377_ssc_1
      | ln_and_242_ssc_1 | ln_and_379_ssc_1 | ln_land_252_lpi_1_dfm_1))) | ln_and_407_ssc_1
      | ln_and_244_ssc_1 | ln_and_246_ssc_1) & ln_nor_9_cse_1;
  assign ln_ln_ln_or_32_nl = (~((~((ln_ln_mux1h_118_psp_1_3 & (~(ln_and_240_ssc_1
      | ln_and_377_ssc_1 | ln_and_242_ssc_1 | ln_and_407_ssc_1 | ln_and_379_ssc_1)))
      | ln_and_244_ssc_1 | ln_and_246_ssc_1 | ln_land_252_lpi_1_dfm_1)) | ln_if_253_acc_cse_11_sva_1))
      | ln_and_248_ssc_1;
  assign ln_ln_ln_or_34_nl = (~((~((ln_ln_mux1h_118_psp_1_2 & (~(ln_and_240_ssc_1
      | ln_and_244_ssc_1 | ln_and_379_ssc_1 | ln_and_246_ssc_1))) | ln_and_377_ssc_1
      | ln_and_242_ssc_1 | ln_and_407_ssc_1 | ln_land_252_lpi_1_dfm_1)) | ln_if_253_acc_cse_11_sva_1))
      | ln_and_248_ssc_1;
  assign ln_ln_ln_or_36_nl = (ln_ln_mux1h_118_psp_1_1 & (~(ln_and_377_ssc_1 | ln_and_407_ssc_1
      | ln_and_244_ssc_1 | ln_land_252_lpi_1_dfm_1))) | ln_and_240_ssc_1 | ln_and_242_ssc_1
      | ln_and_379_ssc_1 | ln_and_246_ssc_1 | ln_and_248_ssc_1 | ln_if_253_acc_cse_11_sva_1;
  assign ln_ln_ln_or_37_nl = (ln_ln_mux1h_118_psp_1_0 & (~(ln_and_240_ssc_1 | ln_and_242_ssc_1
      | ln_and_407_ssc_1 | ln_and_244_ssc_1 | ln_and_246_ssc_1))) | ln_and_377_ssc_1
      | ln_and_379_ssc_1 | ln_land_252_lpi_1_dfm_1 | ln_and_248_ssc_1 | ln_if_253_acc_cse_11_sva_1;
  assign nl_if_4_for_if_if_4_for_if_mul_nl = $signed(({1'b1 , ln_ln_ln_and_4_nl ,
      ln_ln_ln_or_20_nl , ln_ln_ln_or_21_nl , ln_ln_ln_and_5_nl , ln_ln_ln_or_24_nl
      , ln_ln_ln_or_26_nl , ln_ln_ln_or_27_nl , ln_ln_ln_and_6_nl , ln_ln_ln_or_30_nl
      , ln_ln_ln_and_7_nl , ln_ln_ln_or_32_nl , ln_ln_ln_or_34_nl , ln_ln_ln_or_36_nl
      , ln_ln_ln_or_37_nl})) * $signed(conv_u2s_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1));
  assign if_4_for_if_if_4_for_if_mul_nl = nl_if_4_for_if_if_4_for_if_mul_nl[24:0];
  assign nl_if_4_for_if_acc_nl = sum1_1_lpi_1_dfm_1 + (readslicef_25_24_1(if_4_for_if_if_4_for_if_mul_nl));
  assign if_4_for_if_acc_nl = nl_if_4_for_if_acc_nl[23:0];
  assign sum1_1_lpi_1_dfm_2_mx0 = MUX_v_24_2_2(sum1_1_lpi_1_dfm_1, if_4_for_if_acc_nl,
      if_4_for_and_45_itm_1);
  assign ln_1_ln_1_ln_1_and_4_nl = (~(ln_1_land_251_lpi_1_dfm_1 | ln_1_land_252_lpi_1_dfm_1))
      & ln_1_nor_9_cse_1;
  assign ln_1_ln_1_ln_1_or_20_nl = (ln_1_ln_1_mux1h_118_psp_1_12 & ln_1_nor_10_cse_1)
      | ln_1_and_246_ssc_1 | ln_1_land_252_lpi_1_dfm_1 | ln_1_and_248_ssc_1 | ln_1_if_253_acc_cse_11_sva_1;
  assign ln_1_ln_1_ln_1_or_21_nl = (~((~((ln_1_ln_1_mux1h_118_psp_1_11 & ln_1_nor_10_cse_1)
      | ln_1_and_246_ssc_1 | ln_1_land_252_lpi_1_dfm_1)) | ln_1_if_253_acc_cse_11_sva_1))
      | ln_1_and_248_ssc_1;
  assign ln_1_ln_1_ln_1_and_5_nl = ((ln_1_ln_1_mux1h_118_psp_1_10 & (~(ln_1_and_407_ssc_1
      | ln_1_and_244_ssc_1 | ln_1_and_379_ssc_1))) | ln_1_and_240_ssc_1 | ln_1_and_377_ssc_1
      | ln_1_and_242_ssc_1 | ln_1_and_246_ssc_1 | ln_1_land_252_lpi_1_dfm_1) & ln_1_nor_9_cse_1;
  assign ln_1_ln_1_ln_1_or_24_nl = (~((~(ln_1_and_427_itm_1 | ln_1_and_407_ssc_1
      | ln_1_and_246_ssc_1)) | ln_1_and_248_ssc_1)) | ln_1_if_253_acc_cse_11_sva_1;
  assign ln_1_ln_1_ln_1_or_26_nl = (ln_1_ln_1_mux1h_118_psp_1_8 & (~(ln_1_and_240_ssc_1
      | ln_1_and_377_ssc_1 | ln_1_and_242_ssc_1 | ln_1_and_379_ssc_1 | ln_1_and_246_ssc_1
      | ln_1_land_252_lpi_1_dfm_1))) | ln_1_and_407_ssc_1 | ln_1_and_244_ssc_1 |
      ln_1_and_248_ssc_1 | ln_1_if_253_acc_cse_11_sva_1;
  assign ln_1_ln_1_ln_1_or_27_nl = (~((~((ln_1_ln_1_mux1h_118_psp_1_7 & (~(ln_1_and_242_ssc_1
      | ln_1_and_407_ssc_1 | ln_1_land_252_lpi_1_dfm_1))) | ln_1_and_240_ssc_1 |
      ln_1_and_377_ssc_1 | ln_1_and_244_ssc_1 | ln_1_and_379_ssc_1 | ln_1_and_246_ssc_1))
      | ln_1_and_248_ssc_1)) | ln_1_if_253_acc_cse_11_sva_1;
  assign ln_1_ln_1_ln_1_and_6_nl = ((ln_1_ln_1_mux1h_118_psp_1_6 & (~(ln_1_and_377_ssc_1
      | ln_1_and_407_ssc_1 | ln_1_and_379_ssc_1 | ln_1_and_246_ssc_1))) | ln_1_and_240_ssc_1
      | ln_1_and_242_ssc_1 | ln_1_and_244_ssc_1 | ln_1_land_252_lpi_1_dfm_1) & ln_1_nor_9_cse_1;
  assign ln_1_ln_1_ln_1_or_30_nl = (ln_1_ln_1_mux1h_118_psp_1_5 & (~(ln_1_and_240_ssc_1
      | ln_1_and_377_ssc_1 | ln_1_and_242_ssc_1 | ln_1_and_379_ssc_1))) | ln_1_and_407_ssc_1
      | ln_1_and_244_ssc_1 | ln_1_and_246_ssc_1 | ln_1_land_252_lpi_1_dfm_1 | ln_1_and_248_ssc_1
      | ln_1_if_253_acc_cse_11_sva_1;
  assign ln_1_ln_1_ln_1_and_7_nl = ((ln_1_ln_1_mux1h_118_psp_1_4 & (~(ln_1_and_240_ssc_1
      | ln_1_and_377_ssc_1 | ln_1_and_242_ssc_1 | ln_1_and_379_ssc_1 | ln_1_land_252_lpi_1_dfm_1)))
      | ln_1_and_407_ssc_1 | ln_1_and_244_ssc_1 | ln_1_and_246_ssc_1) & ln_1_nor_9_cse_1;
  assign ln_1_ln_1_ln_1_or_32_nl = (~((~((ln_1_ln_1_mux1h_118_psp_1_3 & (~(ln_1_and_240_ssc_1
      | ln_1_and_377_ssc_1 | ln_1_and_242_ssc_1 | ln_1_and_407_ssc_1 | ln_1_and_379_ssc_1)))
      | ln_1_and_244_ssc_1 | ln_1_and_246_ssc_1 | ln_1_land_252_lpi_1_dfm_1)) | ln_1_if_253_acc_cse_11_sva_1))
      | ln_1_and_248_ssc_1;
  assign ln_1_ln_1_ln_1_or_34_nl = (~((~((ln_1_ln_1_mux1h_118_psp_1_2 & (~(ln_1_and_240_ssc_1
      | ln_1_and_244_ssc_1 | ln_1_and_379_ssc_1 | ln_1_and_246_ssc_1))) | ln_1_and_377_ssc_1
      | ln_1_and_242_ssc_1 | ln_1_and_407_ssc_1 | ln_1_land_252_lpi_1_dfm_1)) | ln_1_if_253_acc_cse_11_sva_1))
      | ln_1_and_248_ssc_1;
  assign ln_1_ln_1_ln_1_or_36_nl = (ln_1_ln_1_mux1h_118_psp_1_1 & (~(ln_1_and_377_ssc_1
      | ln_1_and_407_ssc_1 | ln_1_and_244_ssc_1 | ln_1_land_252_lpi_1_dfm_1))) |
      ln_1_and_240_ssc_1 | ln_1_and_242_ssc_1 | ln_1_and_379_ssc_1 | ln_1_and_246_ssc_1
      | ln_1_and_248_ssc_1 | ln_1_if_253_acc_cse_11_sva_1;
  assign ln_1_ln_1_ln_1_or_37_nl = (ln_1_ln_1_mux1h_118_psp_1_0 & (~(ln_1_and_240_ssc_1
      | ln_1_and_242_ssc_1 | ln_1_and_407_ssc_1 | ln_1_and_244_ssc_1 | ln_1_and_246_ssc_1)))
      | ln_1_and_377_ssc_1 | ln_1_and_379_ssc_1 | ln_1_land_252_lpi_1_dfm_1 | ln_1_and_248_ssc_1
      | ln_1_if_253_acc_cse_11_sva_1;
  assign nl_if_4_for_1_if_if_4_for_1_if_mul_nl = $signed(({1'b1 , ln_1_ln_1_ln_1_and_4_nl
      , ln_1_ln_1_ln_1_or_20_nl , ln_1_ln_1_ln_1_or_21_nl , ln_1_ln_1_ln_1_and_5_nl
      , ln_1_ln_1_ln_1_or_24_nl , ln_1_ln_1_ln_1_or_26_nl , ln_1_ln_1_ln_1_or_27_nl
      , ln_1_ln_1_ln_1_and_6_nl , ln_1_ln_1_ln_1_or_30_nl , ln_1_ln_1_ln_1_and_7_nl
      , ln_1_ln_1_ln_1_or_32_nl , ln_1_ln_1_ln_1_or_34_nl , ln_1_ln_1_ln_1_or_36_nl
      , ln_1_ln_1_ln_1_or_37_nl})) * $signed(conv_u2s_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1));
  assign if_4_for_1_if_if_4_for_1_if_mul_nl = nl_if_4_for_1_if_if_4_for_1_if_mul_nl[24:0];
  assign nl_if_4_for_1_if_acc_nl = sum2_1_lpi_1_dfm_1 + (readslicef_25_24_1(if_4_for_1_if_if_4_for_1_if_mul_nl));
  assign if_4_for_1_if_acc_nl = nl_if_4_for_1_if_acc_nl[23:0];
  assign sum2_1_lpi_1_dfm_1_mx0 = MUX_v_24_2_2(sum2_1_lpi_1_dfm_1, if_4_for_1_if_acc_nl,
      operator_24_14_false_AC_TRN_AC_WRAP_1_slc_operator_24_14_false_AC_TRN_AC_WRAP_1_acc_14_svs_1);
  assign if_4_for_and_mdf_sva_1 = exit_if_4_for_lpi_1_dfm_3 & (if_4_for_1_acc_tmp[4]);
  assign nl_operator_24_14_false_AC_TRN_AC_WRAP_1_acc_nl = ({1'b1 , (~ operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)})
      + 15'b000000000000001;
  assign operator_24_14_false_AC_TRN_AC_WRAP_1_acc_nl = nl_operator_24_14_false_AC_TRN_AC_WRAP_1_acc_nl[14:0];
  assign operator_24_14_false_AC_TRN_AC_WRAP_1_acc_itm_14_1 = readslicef_15_1_14(operator_24_14_false_AC_TRN_AC_WRAP_1_acc_nl);
  assign asn_sft_lpi_1_dfm_st_1_mx0 = MUX_v_10_2_2(count_sva, asn_sft_lpi_1_dfm_st_1,
      nor_47_cse);
  assign or_49_nl = or_dcpl_29 | or_dcpl_28;
  assign P2_0_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
      P2_0_1_23_10_sva, or_49_nl);
  assign or_55_nl = or_dcpl_29 | or_dcpl_34;
  assign P2_8_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
      P2_8_1_23_10_sva, or_55_nl);
  assign operator_24_14_false_AC_TRN_AC_WRAP_operator_24_14_false_AC_TRN_AC_WRAP_operator_24_14_false_AC_TRN_AC_WRAP_mux_nl
      = MUX_v_14_16_2(P2_0_1_23_10_sva, P2_1_1_23_10_sva, P2_2_1_23_10_sva, P2_3_1_23_10_sva,
      P2_4_1_23_10_sva, P2_5_1_23_10_sva, P2_6_1_23_10_sva, P2_7_1_23_10_sva, P2_8_1_23_10_sva,
      P2_9_1_23_10_sva, P2_10_1_23_10_sva, P2_11_1_23_10_sva, P2_12_1_23_10_sva,
      P2_13_1_23_10_sva, P2_14_1_23_10_sva, P2_15_1_23_10_sva, {shift_reg_1_sva_2
      , shift_reg_1_sva_1 , shift_reg_1_sva_0 , epsilon_rsci_idat});
  assign nl_operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_operator_24_14_false_AC_TRN_AC_WRAP_operator_24_14_false_AC_TRN_AC_WRAP_mux_nl
      + 14'b00000000000001;
  assign operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1 = nl_operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1[13:0];
  assign or_58_nl = or_dcpl_37 | or_dcpl_28;
  assign P2_1_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
      P2_1_1_23_10_sva, or_58_nl);
  assign or_61_nl = or_dcpl_37 | or_dcpl_34;
  assign P2_9_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
      P2_9_1_23_10_sva, or_61_nl);
  assign or_65_nl = or_dcpl_29 | or_dcpl_44;
  assign P2_2_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
      P2_2_1_23_10_sva, or_65_nl);
  assign or_68_nl = or_dcpl_29 | or_dcpl_47;
  assign P2_10_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
      P2_10_1_23_10_sva, or_68_nl);
  assign or_70_nl = or_dcpl_37 | or_dcpl_44;
  assign P2_3_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
      P2_3_1_23_10_sva, or_70_nl);
  assign or_72_nl = or_dcpl_37 | or_dcpl_47;
  assign P2_11_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
      P2_11_1_23_10_sva, or_72_nl);
  assign or_76_nl = or_dcpl_29 | or_dcpl_55;
  assign P2_12_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
      P2_12_1_23_10_sva, or_76_nl);
  assign or_79_nl = or_dcpl_29 | or_dcpl_58;
  assign P2_4_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
      P2_4_1_23_10_sva, or_79_nl);
  assign or_81_nl = or_dcpl_37 | or_dcpl_55;
  assign P2_13_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
      P2_13_1_23_10_sva, or_81_nl);
  assign or_83_nl = or_dcpl_37 | or_dcpl_58;
  assign P2_5_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
      P2_5_1_23_10_sva, or_83_nl);
  assign or_87_nl = or_dcpl_29 | or_dcpl_66;
  assign P2_14_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
      P2_14_1_23_10_sva, or_87_nl);
  assign or_90_nl = or_dcpl_29 | or_dcpl_69;
  assign P2_6_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
      P2_6_1_23_10_sva, or_90_nl);
  assign or_92_nl = or_dcpl_37 | or_dcpl_66;
  assign P2_15_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
      P2_15_1_23_10_sva, or_92_nl);
  assign or_94_nl = or_dcpl_37 | or_dcpl_69;
  assign P2_7_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
      P2_7_1_23_10_sva, or_94_nl);
  assign or_98_ssc = mux_tmp_4 | or_dcpl_77;
  assign P1_0_1_23_10_sva_dfm_1_mx0_13_12 = MUX_v_2_2_2((operator_24_14_false_AC_TRN_AC_WRAP_1_acc_psp_sva_1[13:12]),
      P1_0_1_23_10_sva_rsp_0, or_98_ssc);
  assign P1_0_1_23_10_sva_dfm_1_mx0_11_0 = MUX_v_12_2_2((operator_24_14_false_AC_TRN_AC_WRAP_1_acc_psp_sva_1[11:0]),
      P1_0_1_23_10_sva_rsp_1, or_98_ssc);
  assign or_102_nl = mux_tmp_4 | or_dcpl_81;
  assign P1_4_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_1_acc_psp_sva_1,
      P1_4_1_23_10_sva, or_102_nl);
  assign operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_nl
      = MUX_v_14_8_2(({P1_0_1_23_10_sva_rsp_0 , P1_0_1_23_10_sva_rsp_1}), P1_1_1_23_10_sva,
      P1_2_1_23_10_sva, P1_3_1_23_10_sva, P1_4_1_23_10_sva, P1_5_1_23_10_sva, P1_6_1_23_10_sva,
      P1_7_1_23_10_sva, {shift_reg_1_sva_1 , shift_reg_1_sva_0 , epsilon_rsci_idat});
  assign nl_operator_24_14_false_AC_TRN_AC_WRAP_1_acc_psp_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_nl
      + 14'b00000000000001;
  assign operator_24_14_false_AC_TRN_AC_WRAP_1_acc_psp_sva_1 = nl_operator_24_14_false_AC_TRN_AC_WRAP_1_acc_psp_sva_1[13:0];
  assign or_104_nl = (~ mux_1310_itm) | or_dcpl_77;
  assign P1_1_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_1_acc_psp_sva_1,
      P1_1_1_23_10_sva, or_104_nl);
  assign or_106_nl = (~ mux_1310_itm) | or_dcpl_81;
  assign P1_5_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_1_acc_psp_sva_1,
      P1_5_1_23_10_sva, or_106_nl);
  assign or_109_nl = mux_tmp_4 | or_dcpl_88;
  assign P1_2_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_1_acc_psp_sva_1,
      P1_2_1_23_10_sva, or_109_nl);
  assign or_112_nl = mux_tmp_4 | or_dcpl_91;
  assign P1_6_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_1_acc_psp_sva_1,
      P1_6_1_23_10_sva, or_112_nl);
  assign or_114_nl = (~ mux_1310_itm) | or_dcpl_88;
  assign P1_3_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_1_acc_psp_sva_1,
      P1_3_1_23_10_sva, or_114_nl);
  assign or_116_nl = (~ mux_1310_itm) | or_dcpl_91;
  assign P1_7_1_23_10_sva_dfm_1_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_1_acc_psp_sva_1,
      P1_7_1_23_10_sva, or_116_nl);
  assign or_135_nl = mux_tmp_11 | or_dcpl_104;
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_mux_3_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_0_2_23_10_sva_mx0, or_135_nl);
  assign or_142_nl = mux_tmp_16 | or_dcpl_104;
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_mux_7_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_1_2_23_10_sva_mx0, or_142_nl);
  assign or_153_nl = mux_tmp_22 | or_dcpl_104;
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_mux_11_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_2_2_23_10_sva_mx0, or_153_nl);
  assign or_159_nl = not_tmp_48 | or_dcpl_104;
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_mux_15_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_3_2_23_10_sva_mx0, or_159_nl);
  assign or_169_nl = mux_tmp_11 | or_dcpl_121;
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_mux_19_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_4_2_23_10_sva_mx0, or_169_nl);
  assign or_177_nl = mux_tmp_16 | or_dcpl_121;
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_mux_23_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_5_2_23_10_sva_mx0, or_177_nl);
  assign or_184_nl = mux_tmp_22 | or_dcpl_121;
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_mux_27_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_6_2_23_10_sva_mx0, or_184_nl);
  assign or_192_nl = not_tmp_48 | or_dcpl_121;
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_mux_31_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_7_2_23_10_sva_mx0, or_192_nl);
  assign or_129_nl = mux_tmp_11 | or_dcpl_98;
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_mux_1_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_8_2_23_10_sva_mx0, or_129_nl);
  assign or_140_nl = mux_tmp_16 | or_dcpl_98;
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_mux_5_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_9_2_23_10_sva_mx0, or_140_nl);
  assign or_151_nl = mux_tmp_22 | or_dcpl_98;
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_mux_9_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_10_2_23_10_sva_mx0, or_151_nl);
  assign or_157_nl = not_tmp_48 | or_dcpl_98;
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_mux_13_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_11_2_23_10_sva_mx0, or_157_nl);
  assign or_162_nl = mux_tmp_11 | or_dcpl_118;
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_mux_17_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_12_2_23_10_sva_mx0, or_162_nl);
  assign or_171_nl = mux_tmp_16 | or_dcpl_118;
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_mux_21_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_13_2_23_10_sva_mx0, or_171_nl);
  assign or_179_nl = mux_tmp_22 | or_dcpl_118;
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_mux_25_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_14_2_23_10_sva_mx0, or_179_nl);
  assign or_189_nl = not_tmp_48 | or_dcpl_118;
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_mux_29_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_15_2_23_10_sva_mx0, or_189_nl);
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_operator_24_14_false_AC_TRN_AC_WRAP_6_operator_24_14_false_AC_TRN_AC_WRAP_6_mux_nl
      = MUX_v_14_16_2(operator_24_14_false_AC_TRN_AC_WRAP_5_mux_3_nl, operator_24_14_false_AC_TRN_AC_WRAP_5_mux_7_nl,
      operator_24_14_false_AC_TRN_AC_WRAP_5_mux_11_nl, operator_24_14_false_AC_TRN_AC_WRAP_5_mux_15_nl,
      operator_24_14_false_AC_TRN_AC_WRAP_5_mux_19_nl, operator_24_14_false_AC_TRN_AC_WRAP_5_mux_23_nl,
      operator_24_14_false_AC_TRN_AC_WRAP_5_mux_27_nl, operator_24_14_false_AC_TRN_AC_WRAP_5_mux_31_nl,
      operator_24_14_false_AC_TRN_AC_WRAP_5_mux_1_nl, operator_24_14_false_AC_TRN_AC_WRAP_5_mux_5_nl,
      operator_24_14_false_AC_TRN_AC_WRAP_5_mux_9_nl, operator_24_14_false_AC_TRN_AC_WRAP_5_mux_13_nl,
      operator_24_14_false_AC_TRN_AC_WRAP_5_mux_17_nl, operator_24_14_false_AC_TRN_AC_WRAP_5_mux_21_nl,
      operator_24_14_false_AC_TRN_AC_WRAP_5_mux_25_nl, operator_24_14_false_AC_TRN_AC_WRAP_5_mux_29_nl,
      {epsilon_rsci_idat , saved_reg_sva_dfm_1_2_mx0 , saved_reg_sva_dfm_1_1_mx0
      , saved_reg_sva_dfm_1_0_mx0});
  assign nl_operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_operator_24_14_false_AC_TRN_AC_WRAP_6_operator_24_14_false_AC_TRN_AC_WRAP_6_mux_nl
      + 14'b00000000000001;
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1 = nl_operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1[13:0];
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_12_nl = (~ operator_24_14_false_AC_TRN_AC_WRAP_2_and_10_cse_sva_1)
      & operator_24_14_false_AC_TRN_AC_WRAP_3_nor_m1c_mx0w0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_or_nl = (operator_24_14_false_AC_TRN_AC_WRAP_2_and_10_cse_sva_1
      & operator_24_14_false_AC_TRN_AC_WRAP_3_nor_m1c_mx0w0) | (operator_24_14_false_AC_TRN_AC_WRAP_2_and_11_cse_sva_1
      & operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_6_mx0w0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_or_1_nl = ((~ or_dcpl_88) & operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_1_mx0w0)
      | ((~ or_dcpl_81) & operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_4_mx0w0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_35_nl = or_dcpl_88 & operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_1_mx0w0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_37_nl = or_dcpl_81 & operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_4_mx0w0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_27_nl = (~ operator_24_14_false_AC_TRN_AC_WRAP_2_and_11_cse_sva_1)
      & operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_6_mx0w0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_operator_24_14_false_AC_TRN_AC_WRAP_3_operator_24_14_false_AC_TRN_AC_WRAP_3_operator_24_14_false_AC_TRN_AC_WRAP_3_mux1h_nl
      = MUX1HOT_v_14_10_2(({P1_0_1_23_10_sva_rsp_0 , P1_0_1_23_10_sva_rsp_1}), operator_24_14_false_AC_TRN_AC_WRAP_2_acc_psp_sva_1,
      P1_1_1_23_10_sva, operator_24_14_false_AC_TRN_AC_WRAP_1_acc_psp_sva_1, P1_2_1_23_10_sva,
      P1_3_1_23_10_sva, P1_4_1_23_10_sva, P1_5_1_23_10_sva, P1_6_1_23_10_sva, P1_7_1_23_10_sva,
      {operator_24_14_false_AC_TRN_AC_WRAP_3_and_12_nl , operator_24_14_false_AC_TRN_AC_WRAP_3_or_nl
      , operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_mx0w0 , operator_24_14_false_AC_TRN_AC_WRAP_3_or_1_nl
      , operator_24_14_false_AC_TRN_AC_WRAP_3_and_35_nl , operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_2_mx0w0
      , operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_3_mx0w0 , operator_24_14_false_AC_TRN_AC_WRAP_3_and_37_nl
      , operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_5_mx0w0 , operator_24_14_false_AC_TRN_AC_WRAP_3_and_27_nl});
  assign nl_operator_24_14_false_AC_TRN_AC_WRAP_3_acc_psp_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_3_operator_24_14_false_AC_TRN_AC_WRAP_3_operator_24_14_false_AC_TRN_AC_WRAP_3_operator_24_14_false_AC_TRN_AC_WRAP_3_mux1h_nl
      + 14'b00000000000001;
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_acc_psp_sva_1 = nl_operator_24_14_false_AC_TRN_AC_WRAP_3_acc_psp_sva_1[13:0];
  assign or_99_tmp = epsilon_rsci_idat | or_dcpl_77;
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_nor_m1c = ~(shift_reg_1_sva_0 | epsilon_rsci_idat
      | saved_reg_sva_dfm_1_2_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_nor_3_cse = ~(epsilon_rsci_idat |
      saved_reg_sva_dfm_1_2_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_m1c_3 = shift_reg_1_sva_0 & operator_24_14_false_AC_TRN_AC_WRAP_2_nor_3_cse;
  assign or_117_tmp = (~ epsilon_rsci_idat) | or_dcpl_91;
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_m1c_6 = shift_reg_1_sva_0 & epsilon_rsci_idat
      & saved_reg_sva_dfm_1_2_mx0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_or_nl = ((~ or_99_tmp) & operator_24_14_false_AC_TRN_AC_WRAP_2_nor_m1c)
      | ((~ or_117_tmp) & operator_24_14_false_AC_TRN_AC_WRAP_2_and_m1c_6);
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_20_nl = or_99_tmp & operator_24_14_false_AC_TRN_AC_WRAP_2_nor_m1c;
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_21_nl = saved_reg_sva_dfm_1_2_mx0
      & (~(shift_reg_1_sva_0 | epsilon_rsci_idat));
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_22_nl = epsilon_rsci_idat & (~(shift_reg_1_sva_0
      | saved_reg_sva_dfm_1_2_mx0));
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_23_nl = epsilon_rsci_idat & saved_reg_sva_dfm_1_2_mx0
      & (~ shift_reg_1_sva_0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_25_nl = shift_reg_1_sva_0 & saved_reg_sva_dfm_1_2_mx0
      & (~ epsilon_rsci_idat);
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_26_nl = shift_reg_1_sva_0 & epsilon_rsci_idat
      & (~ saved_reg_sva_dfm_1_2_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_27_nl = or_117_tmp & operator_24_14_false_AC_TRN_AC_WRAP_2_and_m1c_6;
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_operator_24_14_false_AC_TRN_AC_WRAP_2_operator_24_14_false_AC_TRN_AC_WRAP_2_operator_24_14_false_AC_TRN_AC_WRAP_2_mux1h_nl
      = MUX1HOT_v_14_9_2(operator_24_14_false_AC_TRN_AC_WRAP_1_acc_psp_sva_1, ({P1_0_1_23_10_sva_rsp_0
      , P1_0_1_23_10_sva_rsp_1}), P1_1_1_23_10_sva, P1_2_1_23_10_sva, P1_3_1_23_10_sva,
      P1_4_1_23_10_sva, P1_5_1_23_10_sva, P1_6_1_23_10_sva, P1_7_1_23_10_sva, {operator_24_14_false_AC_TRN_AC_WRAP_2_or_nl
      , operator_24_14_false_AC_TRN_AC_WRAP_2_and_20_nl , operator_24_14_false_AC_TRN_AC_WRAP_2_and_21_nl
      , operator_24_14_false_AC_TRN_AC_WRAP_2_and_22_nl , operator_24_14_false_AC_TRN_AC_WRAP_2_and_23_nl
      , operator_24_14_false_AC_TRN_AC_WRAP_2_and_m1c_3 , operator_24_14_false_AC_TRN_AC_WRAP_2_and_25_nl
      , operator_24_14_false_AC_TRN_AC_WRAP_2_and_26_nl , operator_24_14_false_AC_TRN_AC_WRAP_2_and_27_nl});
  assign nl_operator_24_14_false_AC_TRN_AC_WRAP_2_acc_psp_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_2_operator_24_14_false_AC_TRN_AC_WRAP_2_operator_24_14_false_AC_TRN_AC_WRAP_2_operator_24_14_false_AC_TRN_AC_WRAP_2_mux1h_nl
      + 14'b00000000000001;
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_acc_psp_sva_1 = nl_operator_24_14_false_AC_TRN_AC_WRAP_2_acc_psp_sva_1[13:0];
  assign or_195_nl = or_dcpl_132 | (~(saved_reg_sva_2 & shift_reg_1_sva_1 & shift_reg_1_sva_0));
  assign P2_15_2_23_10_sva_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_15_1_23_10_sva_dfm_1_mx0, or_195_nl);
  assign or_202_nl = mux_tmp_9 | or_dcpl_144;
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_mux_3_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_0_1_23_10_sva_dfm_1_mx0, or_202_nl);
  assign or_206_nl = (~ mux_tmp_9) | or_dcpl_144;
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_mux_7_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_1_1_23_10_sva_dfm_1_mx0, or_206_nl);
  assign or_216_nl = mux_tmp_9 | or_dcpl_154;
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_mux_11_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_2_1_23_10_sva_dfm_1_mx0, or_216_nl);
  assign or_230_nl = (~ mux_tmp_9) | or_dcpl_154;
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_mux_15_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_3_1_23_10_sva_dfm_1_mx0, or_230_nl);
  assign or_246_nl = mux_tmp_9 | or_dcpl_164;
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_mux_19_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_4_1_23_10_sva_dfm_1_mx0, or_246_nl);
  assign or_256_nl = (~ mux_tmp_9) | or_dcpl_164;
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_mux_23_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_5_1_23_10_sva_dfm_1_mx0, or_256_nl);
  assign or_264_nl = mux_tmp_9 | or_dcpl_174;
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_mux_27_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_6_1_23_10_sva_dfm_1_mx0, or_264_nl);
  assign or_269_nl = (~ mux_tmp_9) | or_dcpl_174;
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_mux_31_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_7_1_23_10_sva_dfm_1_mx0, or_269_nl);
  assign or_266_nl = mux_tmp_9 | or_dcpl_170;
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_mux_29_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_8_1_23_10_sva_dfm_1_mx0, or_266_nl);
  assign or_260_nl = (~ mux_tmp_9) | or_dcpl_170;
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_mux_25_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_9_1_23_10_sva_dfm_1_mx0, or_260_nl);
  assign or_252_nl = mux_tmp_9 | or_251_cse;
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_mux_21_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_10_1_23_10_sva_dfm_1_mx0, or_252_nl);
  assign or_237_nl = (~ mux_tmp_9) | or_251_cse;
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_mux_17_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_11_1_23_10_sva_dfm_1_mx0, or_237_nl);
  assign or_224_nl = mux_tmp_9 | or_dcpl_151;
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_mux_13_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_12_1_23_10_sva_dfm_1_mx0, or_224_nl);
  assign or_213_nl = (~ mux_tmp_9) | or_dcpl_151;
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_mux_9_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_13_1_23_10_sva_dfm_1_mx0, or_213_nl);
  assign or_204_nl = mux_tmp_9 | or_dcpl_139;
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_mux_5_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_14_1_23_10_sva_dfm_1_mx0, or_204_nl);
  assign or_197_nl = (~ mux_tmp_9) | or_dcpl_139;
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_mux_1_nl = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_15_1_23_10_sva_dfm_1_mx0, or_197_nl);
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_operator_24_14_false_AC_TRN_AC_WRAP_5_operator_24_14_false_AC_TRN_AC_WRAP_5_mux_nl
      = MUX_v_14_16_2(operator_24_14_false_AC_TRN_AC_WRAP_4_mux_3_nl, operator_24_14_false_AC_TRN_AC_WRAP_4_mux_7_nl,
      operator_24_14_false_AC_TRN_AC_WRAP_4_mux_11_nl, operator_24_14_false_AC_TRN_AC_WRAP_4_mux_15_nl,
      operator_24_14_false_AC_TRN_AC_WRAP_4_mux_19_nl, operator_24_14_false_AC_TRN_AC_WRAP_4_mux_23_nl,
      operator_24_14_false_AC_TRN_AC_WRAP_4_mux_27_nl, operator_24_14_false_AC_TRN_AC_WRAP_4_mux_31_nl,
      operator_24_14_false_AC_TRN_AC_WRAP_4_mux_29_nl, operator_24_14_false_AC_TRN_AC_WRAP_4_mux_25_nl,
      operator_24_14_false_AC_TRN_AC_WRAP_4_mux_21_nl, operator_24_14_false_AC_TRN_AC_WRAP_4_mux_17_nl,
      operator_24_14_false_AC_TRN_AC_WRAP_4_mux_13_nl, operator_24_14_false_AC_TRN_AC_WRAP_4_mux_9_nl,
      operator_24_14_false_AC_TRN_AC_WRAP_4_mux_5_nl, operator_24_14_false_AC_TRN_AC_WRAP_4_mux_1_nl,
      {shift_reg_1_sva_0 , epsilon_rsci_idat , saved_reg_sva_dfm_1_2_mx0 , saved_reg_sva_dfm_1_1_mx0});
  assign nl_operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_5_operator_24_14_false_AC_TRN_AC_WRAP_5_operator_24_14_false_AC_TRN_AC_WRAP_5_mux_nl
      + 14'b00000000000001;
  assign operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1 = nl_operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1[13:0];
  assign or_200_nl = or_dcpl_102 | saved_reg_sva_2 | shift_reg_1_sva_1 | shift_reg_1_sva_0;
  assign P2_0_2_23_10_sva_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_0_1_23_10_sva_dfm_1_mx0, or_200_nl);
  assign mux_1354_nl = MUX_s_1_2_2(or_226_cse, mux_tmp_9, shift_reg_1_sva_1);
  assign or_203_nl = mux_1354_nl | or_dcpl_118;
  assign P2_14_2_23_10_sva_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_14_1_23_10_sva_dfm_1_mx0, or_203_nl);
  assign mux_1355_nl = MUX_s_1_2_2((~ mux_tmp_9), or_222_cse, shift_reg_1_sva_1);
  assign or_205_nl = mux_1355_nl | or_dcpl_104;
  assign P2_1_2_23_10_sva_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_1_1_23_10_sva_dfm_1_mx0, or_205_nl);
  assign mux_1359_nl = MUX_s_1_2_2(mux_tmp_53, epsilon_rsci_idat, shift_reg_1_sva_2);
  assign mux_1363_nl = MUX_s_1_2_2(mux_tmp_57, mux_1359_nl, saved_reg_sva_2);
  assign or_211_nl = mux_1363_nl | or_dcpl_65;
  assign P2_13_2_23_10_sva_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_13_1_23_10_sva_dfm_1_mx0, or_211_nl);
  assign mux_1364_nl = MUX_s_1_2_2(epsilon_rsci_idat, mux_tmp_53, shift_reg_1_sva_2);
  assign mux_1365_nl = MUX_s_1_2_2((~ mux_1364_nl), mux_tmp_57, saved_reg_sva_2);
  assign or_214_nl = mux_1365_nl | or_dcpl_26;
  assign P2_2_2_23_10_sva_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_2_1_23_10_sva_dfm_1_mx0, or_214_nl);
  assign or_222_cse = shift_reg_1_sva_2 | (~ first_sva) | (mux_3_tmp!=2'b00);
  assign or_221_nl = (~ epsilon_rsci_idat) | shift_reg_1_sva_2 | (~ first_sva) |
      (mux_3_tmp!=2'b00);
  assign mux_1368_cse = MUX_s_1_2_2(or_222_cse, or_221_nl, exitL_exit_approx_sva);
  assign or_219_nl = epsilon_rsci_idat | mux_tmp_61;
  assign mux_1367_cse = MUX_s_1_2_2(mux_tmp_61, or_219_nl, exitL_exit_approx_sva);
  assign mux_1369_nl = MUX_s_1_2_2(mux_1368_cse, mux_1367_cse, shift_reg_1_sva_1);
  assign or_223_nl = mux_1369_nl | (~ shift_reg_1_sva_0);
  assign P2_12_2_23_10_sva_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_12_1_23_10_sva_dfm_1_mx0, or_223_nl);
  assign or_226_cse = (~ shift_reg_1_sva_2) | (~ first_sva) | (mux_3_tmp!=2'b00);
  assign and_183_nl = epsilon_rsci_idat & mux_tmp_61;
  assign mux_1372_cse = MUX_s_1_2_2(mux_tmp_61, and_183_nl, exitL_exit_approx_sva);
  assign or_225_nl = epsilon_rsci_idat | (~ shift_reg_1_sva_2) | (~ first_sva) |
      (mux_3_tmp!=2'b00);
  assign mux_1370_nl = MUX_s_1_2_2(or_226_cse, or_225_nl, exitL_exit_approx_sva);
  assign mux_1373_nl = MUX_s_1_2_2((~ mux_1372_cse), mux_1370_nl, shift_reg_1_sva_1);
  assign or_229_nl = mux_1373_nl | shift_reg_1_sva_0;
  assign P2_3_2_23_10_sva_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_3_1_23_10_sva_dfm_1_mx0, or_229_nl);
  assign nor_63_cse = ~((~ shift_reg_1_sva_2) | (~ first_sva) | (mux_3_tmp!=2'b00));
  assign nor_64_nl = ~(epsilon_rsci_idat | (~ shift_reg_1_sva_2) | (~ first_sva)
      | (mux_3_tmp!=2'b00));
  assign mux_1374_nl = MUX_s_1_2_2(nor_63_cse, nor_64_nl, exitL_exit_approx_sva);
  assign mux_1377_nl = MUX_s_1_2_2(mux_1372_cse, mux_1374_nl, shift_reg_1_sva_0);
  assign nand_45_nl = ~(mux_1377_nl & shift_reg_1_sva_1);
  assign P2_11_2_23_10_sva_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_11_1_23_10_sva_dfm_1_mx0, nand_45_nl);
  assign mux_1381_nl = MUX_s_1_2_2(mux_1368_cse, mux_1367_cse, shift_reg_1_sva_0);
  assign or_244_nl = mux_1381_nl | shift_reg_1_sva_1;
  assign P2_4_2_23_10_sva_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_4_1_23_10_sva_dfm_1_mx0, or_244_nl);
  assign or_251_cse = or_dcpl_54 | (~ epsilon_rsci_idat);
  assign or_295_nl = shift_reg_1_sva_1 | (~ shift_reg_1_sva_0) | epsilon_rsci_idat;
  assign mux_1383_cse = MUX_s_1_2_2(or_251_cse, or_295_nl, shift_reg_1_sva_2);
  assign or_247_cse = (~ first_sva) | (mux_3_tmp!=2'b00);
  assign or_249_nl = saved_reg_sva_2 | (~ shift_reg_1_sva_1) | shift_reg_1_sva_0
      | (~ epsilon_rsci_idat);
  assign mux_1384_nl = MUX_s_1_2_2(mux_1383_cse, or_249_nl, or_247_cse);
  assign P2_10_2_23_10_sva_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_10_1_23_10_sva_dfm_1_mx0, mux_1384_nl);
  assign or_293_nl = (~ saved_reg_sva_2) | shift_reg_1_sva_1 | (~ shift_reg_1_sva_0)
      | epsilon_rsci_idat;
  assign mux_1387_nl = MUX_s_1_2_2(mux_1383_cse, or_293_nl, or_247_cse);
  assign P2_5_2_23_10_sva_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_5_1_23_10_sva_dfm_1_mx0, mux_1387_nl);
  assign mux_1388_nl = MUX_s_1_2_2((~ mux_tmp_9), or_222_cse, shift_reg_1_sva_0);
  assign or_258_nl = mux_1388_nl | epsilon_rsci_idat | (~ shift_reg_1_sva_1);
  assign P2_9_2_23_10_sva_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_9_1_23_10_sva_dfm_1_mx0, or_258_nl);
  assign mux_1389_nl = MUX_s_1_2_2(or_226_cse, mux_tmp_9, shift_reg_1_sva_0);
  assign or_262_nl = mux_1389_nl | (~ epsilon_rsci_idat) | shift_reg_1_sva_1;
  assign P2_6_2_23_10_sva_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_6_1_23_10_sva_dfm_1_mx0, or_262_nl);
  assign nand_9_nl = ~(shift_reg_1_sva_1 & (~ mux_tmp_9));
  assign mux_1390_nl = MUX_s_1_2_2(nand_9_nl, or_tmp_12, shift_reg_1_sva_0);
  assign or_265_nl = mux_1390_nl | epsilon_rsci_idat;
  assign P2_8_2_23_10_sva_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_8_1_23_10_sva_dfm_1_mx0, or_265_nl);
  assign or_267_nl = shift_reg_1_sva_1 | (~ mux_tmp_9);
  assign mux_1391_nl = MUX_s_1_2_2(or_tmp_29, or_267_nl, shift_reg_1_sva_0);
  assign or_268_nl = mux_1391_nl | (~ epsilon_rsci_idat);
  assign P2_7_2_23_10_sva_mx0 = MUX_v_14_2_2(operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1,
      P2_7_1_23_10_sva_dfm_1_mx0, or_268_nl);
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_operator_24_14_false_AC_TRN_AC_WRAP_4_operator_24_14_false_AC_TRN_AC_WRAP_4_mux_nl
      = MUX_v_14_16_2(P2_0_1_23_10_sva_dfm_1_mx0, P2_1_1_23_10_sva_dfm_1_mx0, P2_2_1_23_10_sva_dfm_1_mx0,
      P2_3_1_23_10_sva_dfm_1_mx0, P2_4_1_23_10_sva_dfm_1_mx0, P2_5_1_23_10_sva_dfm_1_mx0,
      P2_6_1_23_10_sva_dfm_1_mx0, P2_7_1_23_10_sva_dfm_1_mx0, P2_8_1_23_10_sva_dfm_1_mx0,
      P2_9_1_23_10_sva_dfm_1_mx0, P2_10_1_23_10_sva_dfm_1_mx0, P2_11_1_23_10_sva_dfm_1_mx0,
      P2_12_1_23_10_sva_dfm_1_mx0, P2_13_1_23_10_sva_dfm_1_mx0, P2_14_1_23_10_sva_dfm_1_mx0,
      P2_15_1_23_10_sva_dfm_1_mx0, {shift_reg_1_sva_1 , shift_reg_1_sva_0 , epsilon_rsci_idat
      , saved_reg_sva_dfm_1_2_mx0});
  assign nl_operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_4_operator_24_14_false_AC_TRN_AC_WRAP_4_operator_24_14_false_AC_TRN_AC_WRAP_4_mux_nl
      + 14'b00000000000001;
  assign operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1 = nl_operator_24_14_false_AC_TRN_AC_WRAP_4_acc_psp_sva_1[13:0];
  assign shift_reg_1_sva_0_mx0 = MUX_s_1_2_2(epsilon_rsci_idat, shift_reg_1_sva_0,
      nor_47_cse);
  assign nor_66_nl = ~(reg_skip_ftd | (reg_skip_ftd_1!=2'b00));
  assign skip_sva_dfm_1_0_mx0 = MUX_v_2_2_2(skip_sva_1_1_0_1, reg_skip_ftd_1, nor_66_nl);
  assign saved_reg_sva_dfm_1_2_mx0 = MUX_s_1_2_2(shift_reg_1_sva_2, saved_reg_sva_2,
      or_247_cse);
  assign saved_reg_sva_dfm_1_0_mx0 = MUX_s_1_2_2(shift_reg_1_sva_0, saved_reg_sva_0,
      or_247_cse);
  assign saved_reg_sva_dfm_1_1_mx0 = MUX_s_1_2_2(shift_reg_1_sva_1, saved_reg_sva_1,
      or_247_cse);
  assign nl_skip_sva_1_1_0_1 = reg_skip_ftd_1 + 2'b11;
  assign skip_sva_1_1_0_1 = nl_skip_sva_1_1_0_1[1:0];
  assign or_psp_mx0 = MUX_s_1_2_2(or_324_cse, or_psp, nor_47_cse);
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_0_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_1_0_sva_1
      & (~ saved_reg_sva_dfm_1_2_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_1_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_1_1_sva_1
      & (~ saved_reg_sva_dfm_1_2_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_2_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_1_2_sva_1
      & (~ saved_reg_sva_dfm_1_2_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_3_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_1_3_sva_1
      & (~ saved_reg_sva_dfm_1_2_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_4_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_1_0_sva_1
      & saved_reg_sva_dfm_1_2_mx0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_5_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_1_1_sva_1
      & saved_reg_sva_dfm_1_2_mx0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_6_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_1_2_sva_1
      & saved_reg_sva_dfm_1_2_mx0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_7_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_1_3_sva_1
      & saved_reg_sva_dfm_1_2_mx0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_6_mx0w0 = epsilon_rsci_idat
      & saved_reg_sva_dfm_1_2_mx0 & saved_reg_sva_dfm_1_1_mx0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_6_mx0 = MUX_s_1_2_2(operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_6_mx0w0,
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_6, nor_47_cse);
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_nor_m1c_mx0w0 = ~(epsilon_rsci_idat
      | saved_reg_sva_dfm_1_2_mx0 | saved_reg_sva_dfm_1_1_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_nor_m1c_mx0 = MUX_s_1_2_2(operator_24_14_false_AC_TRN_AC_WRAP_3_nor_m1c_mx0w0,
      operator_24_14_false_AC_TRN_AC_WRAP_3_nor_m1c, nor_47_cse);
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_5_mx0w0 = epsilon_rsci_idat
      & saved_reg_sva_dfm_1_2_mx0 & (~ saved_reg_sva_dfm_1_1_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_5_mx0 = MUX_s_1_2_2(operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_5_mx0w0,
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_5, nor_47_cse);
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_mx0w0 = saved_reg_sva_dfm_1_1_mx0
      & operator_24_14_false_AC_TRN_AC_WRAP_2_nor_3_cse;
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_mx0 = MUX_s_1_2_2(operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_mx0w0,
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c, nor_47_cse);
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_4_mx0w0 = epsilon_rsci_idat
      & saved_reg_sva_dfm_1_1_mx0 & (~ saved_reg_sva_dfm_1_2_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_4_mx0 = MUX_s_1_2_2(operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_4_mx0w0,
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_4, nor_47_cse);
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_1_mx0w0 = saved_reg_sva_dfm_1_2_mx0
      & (~(epsilon_rsci_idat | saved_reg_sva_dfm_1_1_mx0));
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_1_mx0 = MUX_s_1_2_2(operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_1_mx0w0,
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_1, nor_47_cse);
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_3_mx0w0 = epsilon_rsci_idat
      & (~(saved_reg_sva_dfm_1_2_mx0 | saved_reg_sva_dfm_1_1_mx0));
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_3_mx0 = MUX_s_1_2_2(operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_3_mx0w0,
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_3, nor_47_cse);
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_2_mx0w0 = saved_reg_sva_dfm_1_2_mx0
      & saved_reg_sva_dfm_1_1_mx0 & (~ epsilon_rsci_idat);
  assign operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_2_mx0 = MUX_s_1_2_2(operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_2_mx0w0,
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_2, nor_47_cse);
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_11_cse_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_2_and_stg_1_3_sva_1
      & shift_reg_1_sva_0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_10_cse_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_2_nor_3_cse
      & (~ shift_reg_1_sva_0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_9_cse_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_2_and_stg_1_2_sva_1
      & shift_reg_1_sva_0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_8_cse_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_2_and_stg_1_1_sva_1
      & (~ shift_reg_1_sva_0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_7_cse_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_2_and_stg_1_1_sva_1
      & shift_reg_1_sva_0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_6_cse_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_2_and_stg_1_2_sva_1
      & (~ shift_reg_1_sva_0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_4_cse_sva_1 = operator_24_14_false_AC_TRN_AC_WRAP_2_and_stg_1_3_sva_1
      & (~ shift_reg_1_sva_0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_1_0_sva_1 = ~(saved_reg_sva_dfm_1_0_mx0
      | saved_reg_sva_dfm_1_1_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_1_1_sva_1 = saved_reg_sva_dfm_1_0_mx0
      & (~ saved_reg_sva_dfm_1_1_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_1_2_sva_1 = (~ saved_reg_sva_dfm_1_0_mx0)
      & saved_reg_sva_dfm_1_1_mx0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_1_3_sva_1 = saved_reg_sva_dfm_1_0_mx0
      & saved_reg_sva_dfm_1_1_mx0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_stg_1_3_sva_1 = saved_reg_sva_dfm_1_2_mx0
      & epsilon_rsci_idat;
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_stg_1_2_sva_1 = (~ saved_reg_sva_dfm_1_2_mx0)
      & epsilon_rsci_idat;
  assign operator_24_14_false_AC_TRN_AC_WRAP_2_and_stg_1_1_sva_1 = saved_reg_sva_dfm_1_2_mx0
      & (~ epsilon_rsci_idat);
  assign nl_j_1_3_0_sva_2 = conv_u2u_3_4(j_1_3_0_lpi_1_dfm_2_0_1) + 4'b0001;
  assign j_1_3_0_sva_2 = nl_j_1_3_0_sva_2[3:0];
  assign if_4_for_if_4_for_if_4_for_not_3_nl = ~ or_2_tmp;
  assign j_1_3_0_lpi_1_dfm_2_0_1 = MUX_v_3_2_2(3'b000, j_1_3_0_lpi_1_dfm_2_2_0, if_4_for_if_4_for_if_4_for_not_3_nl);
  assign nand_53_ssc = ~((~((~ operator_24_14_false_AC_TRN_AC_WRAP_2_and_10_cse_sva_1)
      & and_7_m1c_1)) & or_2_tmp);
  assign and_76_ssc = operator_24_14_false_AC_TRN_AC_WRAP_2_and_10_cse_sva_1 & and_7_m1c_1;
  assign and_8_ssc = operator_24_14_false_AC_TRN_AC_WRAP_3_nor_m1c_mx0 & or_2_tmp;
  assign P1_0_1_23_10_sva_dfm_3_13_12 = MUX1HOT_v_2_3_2(P1_0_1_23_10_sva_dfm_1_mx0_13_12,
      (operator_24_14_false_AC_TRN_AC_WRAP_2_acc_psp_sva_1[13:12]), (operator_24_14_false_AC_TRN_AC_WRAP_3_acc_psp_sva_1[13:12]),
      {nand_53_ssc , and_76_ssc , and_8_ssc});
  assign P1_0_1_23_10_sva_dfm_3_11_0 = MUX1HOT_v_12_3_2(P1_0_1_23_10_sva_dfm_1_mx0_11_0,
      (operator_24_14_false_AC_TRN_AC_WRAP_2_acc_psp_sva_1[11:0]), (operator_24_14_false_AC_TRN_AC_WRAP_3_acc_psp_sva_1[11:0]),
      {nand_53_ssc , and_76_ssc , and_8_ssc});
  assign nand_55_nl = ~((~((~ operator_24_14_false_AC_TRN_AC_WRAP_2_and_8_cse_sva_1)
      & and_9_m1c_1)) & or_2_tmp);
  assign and_78_nl = operator_24_14_false_AC_TRN_AC_WRAP_2_and_8_cse_sva_1 & and_9_m1c_1;
  assign and_10_nl = operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_mx0 & or_2_tmp;
  assign P1_1_1_23_10_sva_dfm_3 = MUX1HOT_v_14_3_2(P1_1_1_23_10_sva_dfm_1_mx0, operator_24_14_false_AC_TRN_AC_WRAP_2_acc_psp_sva_1,
      operator_24_14_false_AC_TRN_AC_WRAP_3_acc_psp_sva_1, {nand_55_nl , and_78_nl
      , and_10_nl});
  assign nand_57_nl = ~((~((~ operator_24_14_false_AC_TRN_AC_WRAP_2_and_6_cse_sva_1)
      & and_11_m1c_1)) & or_2_tmp);
  assign and_80_nl = operator_24_14_false_AC_TRN_AC_WRAP_2_and_6_cse_sva_1 & and_11_m1c_1;
  assign and_12_nl = operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_1_mx0 & or_2_tmp;
  assign P1_2_1_23_10_sva_dfm_3 = MUX1HOT_v_14_3_2(P1_2_1_23_10_sva_dfm_1_mx0, operator_24_14_false_AC_TRN_AC_WRAP_2_acc_psp_sva_1,
      operator_24_14_false_AC_TRN_AC_WRAP_3_acc_psp_sva_1, {nand_57_nl , and_80_nl
      , and_12_nl});
  assign nand_59_nl = ~((~((~ operator_24_14_false_AC_TRN_AC_WRAP_2_and_4_cse_sva_1)
      & and_13_m1c_1)) & or_2_tmp);
  assign and_82_nl = operator_24_14_false_AC_TRN_AC_WRAP_2_and_4_cse_sva_1 & and_13_m1c_1;
  assign and_14_nl = operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_2_mx0 & or_2_tmp;
  assign P1_3_1_23_10_sva_dfm_3 = MUX1HOT_v_14_3_2(P1_3_1_23_10_sva_dfm_1_mx0, operator_24_14_false_AC_TRN_AC_WRAP_2_acc_psp_sva_1,
      operator_24_14_false_AC_TRN_AC_WRAP_3_acc_psp_sva_1, {nand_59_nl , and_82_nl
      , and_14_nl});
  assign nand_61_nl = ~((~((~ operator_24_14_false_AC_TRN_AC_WRAP_2_and_m1c_3) &
      and_15_m1c_1)) & or_2_tmp);
  assign and_84_nl = operator_24_14_false_AC_TRN_AC_WRAP_2_and_m1c_3 & and_15_m1c_1;
  assign and_16_nl = operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_3_mx0 & or_2_tmp;
  assign P1_4_1_23_10_sva_dfm_3 = MUX1HOT_v_14_3_2(P1_4_1_23_10_sva_dfm_1_mx0, operator_24_14_false_AC_TRN_AC_WRAP_2_acc_psp_sva_1,
      operator_24_14_false_AC_TRN_AC_WRAP_3_acc_psp_sva_1, {nand_61_nl , and_84_nl
      , and_16_nl});
  assign nand_63_nl = ~((~((~ operator_24_14_false_AC_TRN_AC_WRAP_2_and_7_cse_sva_1)
      & and_17_m1c_1)) & or_2_tmp);
  assign and_86_nl = operator_24_14_false_AC_TRN_AC_WRAP_2_and_7_cse_sva_1 & and_17_m1c_1;
  assign and_18_nl = operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_4_mx0 & or_2_tmp;
  assign P1_5_1_23_10_sva_dfm_3 = MUX1HOT_v_14_3_2(P1_5_1_23_10_sva_dfm_1_mx0, operator_24_14_false_AC_TRN_AC_WRAP_2_acc_psp_sva_1,
      operator_24_14_false_AC_TRN_AC_WRAP_3_acc_psp_sva_1, {nand_63_nl , and_86_nl
      , and_18_nl});
  assign nand_65_nl = ~((~((~ operator_24_14_false_AC_TRN_AC_WRAP_2_and_9_cse_sva_1)
      & and_19_m1c_1)) & or_2_tmp);
  assign and_88_nl = operator_24_14_false_AC_TRN_AC_WRAP_2_and_9_cse_sva_1 & and_19_m1c_1;
  assign and_20_nl = operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_5_mx0 & or_2_tmp;
  assign P1_6_1_23_10_sva_dfm_3 = MUX1HOT_v_14_3_2(P1_6_1_23_10_sva_dfm_1_mx0, operator_24_14_false_AC_TRN_AC_WRAP_2_acc_psp_sva_1,
      operator_24_14_false_AC_TRN_AC_WRAP_3_acc_psp_sva_1, {nand_65_nl , and_88_nl
      , and_20_nl});
  assign nand_67_nl = ~((~((~ operator_24_14_false_AC_TRN_AC_WRAP_2_and_11_cse_sva_1)
      & and_21_m1c_1)) & or_2_tmp);
  assign and_90_nl = operator_24_14_false_AC_TRN_AC_WRAP_2_and_11_cse_sva_1 & and_21_m1c_1;
  assign and_22_nl = operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_6_mx0 & or_2_tmp;
  assign P1_7_1_23_10_sva_dfm_3 = MUX1HOT_v_14_3_2(P1_7_1_23_10_sva_dfm_1_mx0, operator_24_14_false_AC_TRN_AC_WRAP_2_acc_psp_sva_1,
      operator_24_14_false_AC_TRN_AC_WRAP_3_acc_psp_sva_1, {nand_67_nl , and_90_nl
      , and_22_nl});
  assign exit_if_4_for_lpi_1_dfm_3 = (j_1_3_0_sva_2[3]) | exit_if_4_for_lpi_1_dfm_4;
  assign nl_if_4_for_1_acc_tmp = conv_u2u_4_5(j_lpi_1_dfm_3_0_1) + 5'b00001;
  assign if_4_for_1_acc_tmp = nl_if_4_for_1_acc_tmp[4:0];
  assign if_4_for_if_4_for_if_4_for_not_20_nl = ~ or_2_tmp;
  assign j_lpi_1_dfm_3_0_1 = MUX_v_4_2_2(4'b0000, j_lpi_1_dfm_1_3_0, if_4_for_if_4_for_if_4_for_not_20_nl);
  assign or_133_tmp = or_dcpl_102 | or_dcpl_100 | shift_reg_1_sva_0;
  assign nor_19_m1c = ~(operator_24_14_false_AC_TRN_AC_WRAP_6_and_26_tmp_1 | (~ or_2_tmp));
  assign and_200_nl = (~ or_133_tmp) & nor_19_m1c;
  assign and_201_nl = or_133_tmp & nor_19_m1c;
  assign and_24_nl = operator_24_14_false_AC_TRN_AC_WRAP_6_and_26_tmp_1 & or_2_tmp;
  assign P2_0_1_23_10_sva_dfm_3 = MUX1HOT_v_14_4_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_0_2_23_10_sva_mx0, operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1,
      P2_0_1_23_10_sva, {and_200_nl , and_201_nl , and_24_nl , (~ or_2_tmp)});
  assign mux_1322_nl = MUX_s_1_2_2(mux_tmp_16, or_tmp_12, shift_reg_1_sva_0);
  assign or_141_tmp = mux_1322_nl | epsilon_rsci_idat;
  assign nor_20_m1c = ~(operator_24_14_false_AC_TRN_AC_WRAP_6_and_24_tmp_1 | (~ or_2_tmp));
  assign and_202_nl = (~ or_141_tmp) & nor_20_m1c;
  assign and_203_nl = or_141_tmp & nor_20_m1c;
  assign and_26_nl = operator_24_14_false_AC_TRN_AC_WRAP_6_and_24_tmp_1 & or_2_tmp;
  assign P2_1_1_23_10_sva_dfm_3 = MUX1HOT_v_14_4_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_1_2_23_10_sva_mx0, operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1,
      P2_1_1_23_10_sva, {and_202_nl , and_203_nl , and_26_nl , (~ or_2_tmp)});
  assign mux_1330_nl = MUX_s_1_2_2(mux_tmp_9, mux_tmp_24, shift_reg_1_sva_1);
  assign mux_1331_nl = MUX_s_1_2_2((~ mux_1330_nl), mux_tmp_23, saved_reg_sva_1);
  assign or_152_tmp = mux_1331_nl | or_dcpl_104;
  assign nor_21_m1c = ~(operator_24_14_false_AC_TRN_AC_WRAP_6_and_22_tmp_1 | (~ or_2_tmp));
  assign and_204_nl = (~ or_152_tmp) & nor_21_m1c;
  assign and_205_nl = or_152_tmp & nor_21_m1c;
  assign and_28_nl = operator_24_14_false_AC_TRN_AC_WRAP_6_and_22_tmp_1 & or_2_tmp;
  assign P2_2_1_23_10_sva_dfm_3 = MUX1HOT_v_14_4_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_2_2_23_10_sva_mx0, operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1,
      P2_2_1_23_10_sva, {and_204_nl , and_205_nl , and_28_nl , (~ or_2_tmp)});
  assign mux_1337_nl = MUX_s_1_2_2(not_tmp_48, or_tmp_19, shift_reg_1_sva_0);
  assign or_158_tmp = mux_1337_nl | epsilon_rsci_idat;
  assign nor_22_m1c = ~(operator_24_14_false_AC_TRN_AC_WRAP_6_and_20_tmp_1 | (~ or_2_tmp));
  assign and_206_nl = (~ or_158_tmp) & nor_22_m1c;
  assign and_207_nl = or_158_tmp & nor_22_m1c;
  assign and_30_nl = operator_24_14_false_AC_TRN_AC_WRAP_6_and_20_tmp_1 & or_2_tmp;
  assign P2_3_1_23_10_sva_dfm_3 = MUX1HOT_v_14_4_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_3_2_23_10_sva_mx0, operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1,
      P2_3_1_23_10_sva, {and_206_nl , and_207_nl , and_30_nl , (~ or_2_tmp)});
  assign mux_1340_nl = MUX_s_1_2_2((~ epsilon_rsci_idat), epsilon_rsci_idat, shift_reg_1_sva_2);
  assign or_166_nl = shift_reg_1_sva_1 | mux_1340_nl;
  assign or_165_nl = or_dcpl_100 | (~ epsilon_rsci_idat);
  assign mux_1341_nl = MUX_s_1_2_2(or_166_nl, or_165_nl, or_247_cse);
  assign or_167_tmp = mux_1341_nl | shift_reg_1_sva_0;
  assign nor_23_m1c = ~(operator_24_14_false_AC_TRN_AC_WRAP_6_and_18_tmp_1 | (~ or_2_tmp));
  assign and_208_nl = (~ or_167_tmp) & nor_23_m1c;
  assign and_209_nl = or_167_tmp & nor_23_m1c;
  assign and_32_nl = operator_24_14_false_AC_TRN_AC_WRAP_6_and_18_tmp_1 & or_2_tmp;
  assign P2_4_1_23_10_sva_dfm_3 = MUX1HOT_v_14_4_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_4_2_23_10_sva_mx0, operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1,
      P2_4_1_23_10_sva, {and_208_nl , and_209_nl , and_32_nl , (~ or_2_tmp)});
  assign or_176_nl = shift_reg_1_sva_2 | (~ and_tmp);
  assign or_175_nl = saved_reg_sva_2 | (~(saved_reg_sva_1 & epsilon_rsci_idat));
  assign mux_1345_nl = MUX_s_1_2_2(or_176_nl, or_175_nl, or_247_cse);
  assign or_173_nl = (~ first_sva) | (mux_3_tmp!=2'b00) | (~ shift_reg_1_sva_2) |
      shift_reg_1_sva_1 | epsilon_rsci_idat;
  assign mux_1346_tmp = MUX_s_1_2_2(mux_1345_nl, or_173_nl, shift_reg_1_sva_0);
  assign nor_24_m1c = ~(operator_24_14_false_AC_TRN_AC_WRAP_6_and_16_tmp_1 | (~ or_2_tmp));
  assign and_210_nl = (~ mux_1346_tmp) & nor_24_m1c;
  assign and_211_nl = mux_1346_tmp & nor_24_m1c;
  assign and_34_nl = operator_24_14_false_AC_TRN_AC_WRAP_6_and_16_tmp_1 & or_2_tmp;
  assign P2_5_1_23_10_sva_dfm_3 = MUX1HOT_v_14_4_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_5_2_23_10_sva_mx0, operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1,
      P2_5_1_23_10_sva, {and_210_nl , and_211_nl , and_34_nl , (~ or_2_tmp)});
  assign mux_1349_nl = MUX_s_1_2_2(epsilon_rsci_idat, (~ epsilon_rsci_idat), shift_reg_1_sva_1);
  assign nand_4_nl = ~(shift_reg_1_sva_2 & mux_1349_nl);
  assign or_182_nl = or_tmp_21 | (~ epsilon_rsci_idat);
  assign mux_1350_nl = MUX_s_1_2_2(nand_4_nl, or_182_nl, or_247_cse);
  assign or_183_tmp = mux_1350_nl | shift_reg_1_sva_0;
  assign nor_25_m1c = ~(operator_24_14_false_AC_TRN_AC_WRAP_6_and_14_tmp_1 | (~ or_2_tmp));
  assign and_212_nl = (~ or_183_tmp) & nor_25_m1c;
  assign and_213_nl = or_183_tmp & nor_25_m1c;
  assign and_36_nl = operator_24_14_false_AC_TRN_AC_WRAP_6_and_14_tmp_1 & or_2_tmp;
  assign P2_6_1_23_10_sva_dfm_3 = MUX1HOT_v_14_4_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_6_2_23_10_sva_mx0, operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1,
      P2_6_1_23_10_sva, {and_212_nl , and_213_nl , and_36_nl , (~ or_2_tmp)});
  assign mux_1352_nl = MUX_s_1_2_2(epsilon_rsci_idat, (~ epsilon_rsci_idat), shift_reg_1_sva_0);
  assign nand_5_nl = ~(shift_reg_1_sva_2 & shift_reg_1_sva_1 & mux_1352_nl);
  assign or_191_nl = shift_reg_1_sva_0 | (~(nor_tmp_5 & epsilon_rsci_idat));
  assign mux_1353_tmp = MUX_s_1_2_2(nand_5_nl, or_191_nl, or_247_cse);
  assign nor_26_m1c = ~(operator_24_14_false_AC_TRN_AC_WRAP_6_and_12_tmp_1 | (~ or_2_tmp));
  assign and_214_nl = (~ mux_1353_tmp) & nor_26_m1c;
  assign and_215_nl = mux_1353_tmp & nor_26_m1c;
  assign and_38_nl = operator_24_14_false_AC_TRN_AC_WRAP_6_and_12_tmp_1 & or_2_tmp;
  assign P2_7_1_23_10_sva_dfm_3 = MUX1HOT_v_14_4_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_7_2_23_10_sva_mx0, operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1,
      P2_7_1_23_10_sva, {and_214_nl , and_215_nl , and_38_nl , (~ or_2_tmp)});
  assign mux_1312_nl = MUX_s_1_2_2((~ epsilon_rsci_idat), epsilon_rsci_idat, shift_reg_1_sva_0);
  assign or_122_nl = shift_reg_1_sva_2 | shift_reg_1_sva_1 | mux_1312_nl;
  assign or_120_nl = (~ shift_reg_1_sva_0) | saved_reg_sva_2 | saved_reg_sva_1 |
      epsilon_rsci_idat;
  assign mux_1313_tmp = MUX_s_1_2_2(or_122_nl, or_120_nl, or_247_cse);
  assign nor_27_m1c = ~(operator_24_14_false_AC_TRN_AC_WRAP_6_and_13_tmp_1 | (~ or_2_tmp));
  assign and_216_nl = (~ mux_1313_tmp) & nor_27_m1c;
  assign and_217_nl = mux_1313_tmp & nor_27_m1c;
  assign and_40_nl = operator_24_14_false_AC_TRN_AC_WRAP_6_and_13_tmp_1 & or_2_tmp;
  assign P2_8_1_23_10_sva_dfm_3 = MUX1HOT_v_14_4_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_8_2_23_10_sva_mx0, operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1,
      P2_8_1_23_10_sva, {and_216_nl , and_217_nl , and_40_nl , (~ or_2_tmp)});
  assign mux_1318_nl = MUX_s_1_2_2((~ epsilon_rsci_idat), epsilon_rsci_idat, shift_reg_1_sva_1);
  assign nor_61_nl = ~(shift_reg_1_sva_2 | mux_1318_nl);
  assign nor_62_nl = ~(saved_reg_sva_2 | (~ saved_reg_sva_1) | epsilon_rsci_idat);
  assign mux_1319_nl = MUX_s_1_2_2(nor_61_nl, nor_62_nl, or_247_cse);
  assign nand_37_tmp = ~(mux_1319_nl & shift_reg_1_sva_0);
  assign nor_28_m1c = ~(operator_24_14_false_AC_TRN_AC_WRAP_6_and_15_tmp_1 | (~ or_2_tmp));
  assign and_218_nl = (~ nand_37_tmp) & nor_28_m1c;
  assign and_219_nl = nand_37_tmp & nor_28_m1c;
  assign and_42_nl = operator_24_14_false_AC_TRN_AC_WRAP_6_and_15_tmp_1 & or_2_tmp;
  assign P2_9_1_23_10_sva_dfm_3 = MUX1HOT_v_14_4_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_9_2_23_10_sva_mx0, operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1,
      P2_9_1_23_10_sva, {and_218_nl , and_219_nl , and_42_nl , (~ or_2_tmp)});
  assign or_149_nl = (~ first_sva) | (mux_3_tmp!=2'b00) | shift_reg_1_sva_2 | (~
      and_tmp);
  assign or_147_nl = (~ shift_reg_1_sva_2) | shift_reg_1_sva_1 | epsilon_rsci_idat;
  assign or_145_nl = or_tmp_21 | epsilon_rsci_idat;
  assign mux_1324_nl = MUX_s_1_2_2(or_147_nl, or_145_nl, or_247_cse);
  assign mux_1325_tmp = MUX_s_1_2_2(or_149_nl, mux_1324_nl, shift_reg_1_sva_0);
  assign nor_29_m1c = ~(operator_24_14_false_AC_TRN_AC_WRAP_6_and_17_tmp_1 | (~ or_2_tmp));
  assign and_220_nl = (~ mux_1325_tmp) & nor_29_m1c;
  assign and_221_nl = mux_1325_tmp & nor_29_m1c;
  assign and_44_nl = operator_24_14_false_AC_TRN_AC_WRAP_6_and_17_tmp_1 & or_2_tmp;
  assign P2_10_1_23_10_sva_dfm_3 = MUX1HOT_v_14_4_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_10_2_23_10_sva_mx0, operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1,
      P2_10_1_23_10_sva, {and_220_nl , and_221_nl , and_44_nl , (~ or_2_tmp)});
  assign mux_1333_nl = MUX_s_1_2_2(epsilon_rsci_idat, (~ epsilon_rsci_idat), shift_reg_1_sva_2);
  assign and_197_nl = shift_reg_1_sva_1 & mux_1333_nl;
  assign and_198_nl = nor_tmp_5 & (~ epsilon_rsci_idat);
  assign mux_1334_nl = MUX_s_1_2_2(and_197_nl, and_198_nl, or_247_cse);
  assign nand_38_tmp = ~(mux_1334_nl & shift_reg_1_sva_0);
  assign nor_30_m1c = ~(operator_24_14_false_AC_TRN_AC_WRAP_6_and_19_tmp_1 | (~ or_2_tmp));
  assign and_222_nl = (~ nand_38_tmp) & nor_30_m1c;
  assign and_223_nl = nand_38_tmp & nor_30_m1c;
  assign and_46_nl = operator_24_14_false_AC_TRN_AC_WRAP_6_and_19_tmp_1 & or_2_tmp;
  assign P2_11_1_23_10_sva_dfm_3 = MUX1HOT_v_14_4_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_11_2_23_10_sva_mx0, operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1,
      P2_11_1_23_10_sva, {and_222_nl , and_223_nl , and_46_nl , (~ or_2_tmp)});
  assign mux_1338_nl = MUX_s_1_2_2(or_tmp_27, mux_tmp_11, shift_reg_1_sva_0);
  assign or_160_tmp = mux_1338_nl | (~ epsilon_rsci_idat);
  assign nor_31_m1c = ~(operator_24_14_false_AC_TRN_AC_WRAP_6_and_21_tmp_1 | (~ or_2_tmp));
  assign and_224_nl = (~ or_160_tmp) & nor_31_m1c;
  assign and_225_nl = or_160_tmp & nor_31_m1c;
  assign and_48_nl = operator_24_14_false_AC_TRN_AC_WRAP_6_and_21_tmp_1 & or_2_tmp;
  assign P2_12_1_23_10_sva_dfm_3 = MUX1HOT_v_14_4_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_12_2_23_10_sva_mx0, operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1,
      P2_12_1_23_10_sva, {and_224_nl , and_225_nl , and_48_nl , (~ or_2_tmp)});
  assign mux_1342_nl = MUX_s_1_2_2(mux_tmp_24, mux_tmp_9, shift_reg_1_sva_1);
  assign mux_1343_nl = MUX_s_1_2_2(mux_tmp_23, mux_1342_nl, saved_reg_sva_1);
  assign or_170_tmp = mux_1343_nl | or_dcpl_118;
  assign nor_32_m1c = ~(operator_24_14_false_AC_TRN_AC_WRAP_6_and_23_tmp_1 | (~ or_2_tmp));
  assign and_226_nl = (~ or_170_tmp) & nor_32_m1c;
  assign and_227_nl = or_170_tmp & nor_32_m1c;
  assign and_50_nl = operator_24_14_false_AC_TRN_AC_WRAP_6_and_23_tmp_1 & or_2_tmp;
  assign P2_13_1_23_10_sva_dfm_3 = MUX1HOT_v_14_4_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_13_2_23_10_sva_mx0, operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1,
      P2_13_1_23_10_sva, {and_226_nl , and_227_nl , and_50_nl , (~ or_2_tmp)});
  assign mux_1347_nl = MUX_s_1_2_2(or_tmp_29, mux_tmp_22, shift_reg_1_sva_0);
  assign or_178_tmp = mux_1347_nl | (~ epsilon_rsci_idat);
  assign nor_33_m1c = ~(operator_24_14_false_AC_TRN_AC_WRAP_6_and_25_tmp_1 | (~ or_2_tmp));
  assign and_228_nl = (~ or_178_tmp) & nor_33_m1c;
  assign and_229_nl = or_178_tmp & nor_33_m1c;
  assign and_52_nl = operator_24_14_false_AC_TRN_AC_WRAP_6_and_25_tmp_1 & or_2_tmp;
  assign P2_14_1_23_10_sva_dfm_3 = MUX1HOT_v_14_4_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_14_2_23_10_sva_mx0, operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1,
      P2_14_1_23_10_sva, {and_228_nl , and_229_nl , and_52_nl , (~ or_2_tmp)});
  assign or_188_tmp = or_dcpl_132 | (~(saved_reg_sva_2 & saved_reg_sva_1 & shift_reg_1_sva_0));
  assign nor_34_m1c = ~(operator_24_14_false_AC_TRN_AC_WRAP_6_and_27_tmp_1 | (~ or_2_tmp));
  assign and_230_nl = (~ or_188_tmp) & nor_34_m1c;
  assign and_231_nl = or_188_tmp & nor_34_m1c;
  assign and_54_nl = operator_24_14_false_AC_TRN_AC_WRAP_6_and_27_tmp_1 & or_2_tmp;
  assign P2_15_1_23_10_sva_dfm_3 = MUX1HOT_v_14_4_2(operator_24_14_false_AC_TRN_AC_WRAP_5_acc_psp_sva_1,
      P2_15_2_23_10_sva_mx0, operator_24_14_false_AC_TRN_AC_WRAP_6_acc_psp_sva_1,
      P2_15_1_23_10_sva, {and_230_nl , and_231_nl , and_54_nl , (~ or_2_tmp)});
  assign exit_if_4_for_lpi_1_dfm_4 = exit_if_4_for_lpi_1_dfm_2 & (~ or_2_tmp);
  assign or_288_nl = or_dcpl_188 | or_dcpl_185 | (if_4_for_mux_50_tmp[9:5]!=5'b11111);
  assign exit_if_4_for_lpi_1_dfm_mx0 = MUX_s_1_2_2(exit_if_4_for_lpi_1_dfm_4, exit_if_4_for_lpi_1_dfm,
      or_288_nl);
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_27_tmp_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_7_sva_1
      & shift_reg_1_sva_0_mx0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_25_tmp_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_6_sva_1
      & shift_reg_1_sva_0_mx0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_23_tmp_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_5_sva_1
      & shift_reg_1_sva_0_mx0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_21_tmp_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_4_sva_1
      & shift_reg_1_sva_0_mx0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_19_tmp_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_3_sva_1
      & shift_reg_1_sva_0_mx0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_17_tmp_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_2_sva_1
      & shift_reg_1_sva_0_mx0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_15_tmp_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_1_sva_1
      & shift_reg_1_sva_0_mx0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_13_tmp_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_0_sva_1
      & shift_reg_1_sva_0_mx0;
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_12_tmp_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_7_sva_1
      & (~ shift_reg_1_sva_0_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_14_tmp_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_6_sva_1
      & (~ shift_reg_1_sva_0_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_16_tmp_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_5_sva_1
      & (~ shift_reg_1_sva_0_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_18_tmp_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_4_sva_1
      & (~ shift_reg_1_sva_0_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_20_tmp_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_3_sva_1
      & (~ shift_reg_1_sva_0_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_22_tmp_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_2_sva_1
      & (~ shift_reg_1_sva_0_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_24_tmp_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_1_sva_1
      & (~ shift_reg_1_sva_0_mx0);
  assign operator_24_14_false_AC_TRN_AC_WRAP_6_and_26_tmp_1 = operator_24_14_false_AC_TRN_AC_WRAP_6_and_stg_2_0_sva_1
      & (~ shift_reg_1_sva_0_mx0);
  assign and_21_m1c_1 = ~(operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_6_mx0 | (~
      or_2_tmp));
  assign and_19_m1c_1 = ~(operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_5_mx0 | (~
      or_2_tmp));
  assign and_17_m1c_1 = ~(operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_4_mx0 | (~
      or_2_tmp));
  assign and_15_m1c_1 = ~(operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_3_mx0 | (~
      or_2_tmp));
  assign and_13_m1c_1 = ~(operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_2_mx0 | (~
      or_2_tmp));
  assign and_11_m1c_1 = ~(operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_1_mx0 | (~
      or_2_tmp));
  assign and_9_m1c_1 = ~(operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_mx0 | (~ or_2_tmp));
  assign and_7_m1c_1 = ~(operator_24_14_false_AC_TRN_AC_WRAP_3_nor_m1c_mx0 | (~ or_2_tmp));
  assign exitL_exit_if_4_for_2_lpi_1_dfm_1 = if_4_for_and_mdf_sva_1 | nand_tmp;
  assign nand_tmp = ~((asn_sft_lpi_1_dfm_st_1_mx0==10'b1111111111));
  assign or_2_tmp = exitL_exit_if_4_for_2_lpi_1_dfm | exitL_exit_approx_sva;
  assign and_55_cse_1 = exit_if_4_for_lpi_1_dfm_mx0 & (~ nand_tmp);
  assign nor_cse_1 = ~(exit_if_4_for_lpi_1_dfm_mx0 | nand_tmp);
  assign and_91_tmp_1 = if_4_for_and_mdf_sva_1 & (~ nand_tmp);
  assign ln_nor_33_cse_1 = ~((~(ln_land_3_lpi_1_dfm_1 | ln_land_4_lpi_1_dfm_1 | ln_and_2_ssc_1))
      | ln_land_6_lpi_1_dfm_1);
  assign ln_land_17_lpi_1_dfm_1 = ln_if_16_acc_itm_12_1 & (~ ln_if_17_acc_itm_14_1);
  assign ln_land_18_lpi_1_dfm_1 = ln_if_17_acc_itm_14_1 & (~ ln_if_18_acc_itm_14_1);
  assign ln_land_19_lpi_1_dfm_1 = ln_if_18_acc_itm_14_1 & (~ ln_if_19_acc_itm_13_1);
  assign ln_land_20_lpi_1_dfm_1 = ln_if_19_acc_itm_13_1 & (~ ln_if_20_acc_itm_14_1);
  assign ln_land_21_lpi_1_dfm_1 = ln_if_20_acc_itm_14_1 & (~ ln_if_21_acc_itm_12_1);
  assign ln_land_22_lpi_1_dfm_1 = ln_if_21_acc_itm_12_1 & (~ ln_if_22_acc_itm_14_1);
  assign ln_land_23_lpi_1_dfm_1 = ln_if_22_acc_itm_14_1 & (~ ln_if_23_acc_itm_13_1);
  assign ln_land_24_lpi_1_dfm_1 = ln_if_23_acc_itm_13_1 & (~ ln_if_24_acc_itm_14_1);
  assign ln_land_25_lpi_1_dfm_1 = ln_if_24_acc_itm_14_1 & (~ ln_if_25_acc_itm_14_1);
  assign ln_land_26_lpi_1_dfm_1 = ln_if_25_acc_itm_14_1 & (~ ln_if_26_acc_itm_12_1);
  assign ln_land_27_lpi_1_dfm_1 = ln_if_26_acc_itm_12_1 & (~ ln_if_27_acc_itm_14_1);
  assign ln_land_28_lpi_1_dfm_1 = ln_if_27_acc_itm_14_1 & (~ ln_if_28_acc_itm_13_1);
  assign ln_land_29_lpi_1_dfm_1 = ln_if_28_acc_itm_13_1 & (~ ln_if_29_acc_itm_14_1);
  assign ln_land_30_lpi_1_dfm_1 = ln_if_29_acc_itm_14_1 & (~ ln_if_30_acc_itm_11_1);
  assign ln_land_31_lpi_1_dfm_1 = ln_if_30_acc_itm_11_1 & (~ ln_if_31_acc_itm_14_1);
  assign ln_land_32_lpi_1_dfm_1 = ln_if_31_acc_itm_14_1 & (~ ln_if_32_acc_itm_14_1);
  assign ln_land_33_lpi_1_dfm_1 = ln_if_32_acc_itm_14_1 & (~ ln_if_33_acc_itm_13_1);
  assign ln_land_34_lpi_1_dfm_1 = ln_if_33_acc_itm_13_1 & (~ ln_if_34_acc_itm_14_1);
  assign ln_land_35_lpi_1_dfm_1 = ln_if_34_acc_itm_14_1 & (~ ln_if_35_acc_itm_11_1);
  assign ln_land_36_lpi_1_dfm_1 = ln_if_35_acc_itm_11_1 & (~ ln_if_36_acc_itm_14_1);
  assign ln_land_37_lpi_1_dfm_1 = ln_if_36_acc_itm_14_1 & (~ ln_if_37_acc_itm_13_1);
  assign ln_land_38_lpi_1_dfm_1 = ln_if_37_acc_itm_13_1 & (~ ln_if_38_acc_itm_14_1);
  assign ln_land_39_lpi_1_dfm_1 = ln_if_38_acc_itm_14_1 & (~ ln_if_39_acc_itm_14_1);
  assign ln_land_40_lpi_1_dfm_1 = ln_if_39_acc_itm_14_1 & (~ ln_if_40_acc_itm_11_1);
  assign ln_land_41_lpi_1_dfm_1 = ln_if_40_acc_itm_11_1 & (~ ln_if_41_acc_itm_14_1);
  assign ln_land_42_lpi_1_dfm_1 = ln_if_41_acc_itm_14_1 & (~ ln_if_42_acc_itm_13_1);
  assign ln_land_43_lpi_1_dfm_1 = ln_if_42_acc_itm_13_1 & (~ ln_if_43_acc_itm_14_1);
  assign ln_land_44_lpi_1_dfm_1 = ln_if_43_acc_itm_14_1 & (~ ln_if_44_acc_itm_12_1);
  assign ln_land_45_lpi_1_dfm_1 = ln_if_44_acc_itm_12_1 & (~ ln_if_45_acc_itm_14_1);
  assign ln_land_46_lpi_1_dfm_1 = ln_if_45_acc_itm_14_1 & (~ ln_if_46_acc_itm_14_1);
  assign ln_land_47_lpi_1_dfm_1 = ln_if_46_acc_itm_14_1 & (~ ln_if_47_acc_itm_13_1);
  assign ln_land_48_lpi_1_dfm_1 = ln_if_47_acc_itm_13_1 & (~ ln_if_48_acc_itm_14_1);
  assign ln_land_49_lpi_1_dfm_1 = ln_if_48_acc_itm_14_1 & (~ ln_if_49_acc_itm_12_1);
  assign ln_if_50_ln_if_50_and_seb_1 = ln_if_49_acc_itm_12_1 & (~ ln_if_50_acc_itm_14_1);
  assign ln_land_51_lpi_1_dfm_1 = ln_if_50_acc_itm_14_1 & (~ ln_if_51_acc_itm_13_1);
  assign ln_land_52_lpi_1_dfm_1 = ln_if_51_acc_itm_13_1 & (~ ln_if_52_acc_itm_14_1);
  assign ln_land_77_lpi_1_dfm_1 = ln_if_76_acc_itm_14_1 & (~ ln_if_77_acc_itm_12_1);
  assign ln_land_78_lpi_1_dfm_1 = ln_if_77_acc_itm_12_1 & (~ ln_if_78_acc_itm_14_1);
  assign ln_land_79_lpi_1_dfm_1 = ln_if_78_acc_itm_14_1 & (~ ln_if_79_acc_itm_13_1);
  assign ln_land_80_lpi_1_dfm_1 = ln_if_79_acc_itm_13_1 & (~ ln_if_80_acc_itm_14_1);
  assign ln_land_81_lpi_1_dfm_1 = ln_if_80_acc_itm_14_1 & (~ ln_if_81_acc_itm_14_1);
  assign ln_land_82_lpi_1_dfm_1 = ln_if_81_acc_itm_14_1 & (~ ln_if_82_acc_itm_12_1);
  assign ln_land_83_lpi_1_dfm_1 = ln_if_82_acc_itm_12_1 & (~ ln_if_83_acc_itm_14_1);
  assign ln_land_84_lpi_1_dfm_1 = ln_if_83_acc_itm_14_1 & (~ ln_if_84_acc_itm_13_1);
  assign ln_land_85_lpi_1_dfm_1 = ln_if_84_acc_itm_13_1 & (~ ln_if_85_acc_itm_14_1);
  assign ln_land_86_lpi_1_dfm_1 = ln_if_85_acc_itm_14_1 & (~ ln_if_86_acc_itm_11_1);
  assign ln_land_87_lpi_1_dfm_1 = ln_if_86_acc_itm_11_1 & (~ ln_if_87_acc_itm_14_1);
  assign ln_land_88_lpi_1_dfm_1 = ln_if_87_acc_itm_14_1 & (~ ln_if_88_acc_itm_14_1);
  assign ln_land_89_lpi_1_dfm_1 = ln_if_88_acc_itm_14_1 & (~ ln_if_89_acc_itm_13_1);
  assign ln_land_90_lpi_1_dfm_1 = ln_if_89_acc_itm_13_1 & (~ ln_if_90_acc_itm_14_1);
  assign ln_land_91_lpi_1_dfm_1 = ln_if_90_acc_itm_14_1 & (~ ln_if_91_acc_itm_11_1);
  assign ln_land_92_lpi_1_dfm_1 = ln_if_91_acc_itm_11_1 & (~ ln_if_92_acc_itm_14_1);
  assign ln_land_93_lpi_1_dfm_1 = ln_if_92_acc_itm_14_1 & (~ ln_if_93_acc_itm_13_1);
  assign ln_land_94_lpi_1_dfm_1 = ln_if_93_acc_itm_13_1 & (~ ln_if_94_acc_itm_14_1);
  assign ln_land_95_lpi_1_dfm_1 = ln_if_94_acc_itm_14_1 & (~ ln_if_95_acc_itm_14_1);
  assign ln_land_96_lpi_1_dfm_1 = ln_if_95_acc_itm_14_1 & (~ ln_if_96_acc_itm_11_1);
  assign ln_land_97_lpi_1_dfm_1 = ln_if_96_acc_itm_11_1 & (~ ln_if_97_acc_itm_14_1);
  assign ln_land_114_lpi_1_dfm_1 = ln_if_113_acc_itm_14_1 & (~ ln_if_114_acc_itm_10_1);
  assign ln_land_115_lpi_1_dfm_1 = ln_if_114_acc_itm_10_1 & (~ ln_if_115_acc_itm_14_1);
  assign ln_land_116_lpi_1_dfm_1 = ln_if_115_acc_itm_14_1 & (~ ln_if_116_acc_itm_14_1);
  assign ln_land_117_lpi_1_dfm_1 = ln_if_116_acc_itm_14_1 & (~ ln_if_117_acc_itm_13_1);
  assign ln_land_118_lpi_1_dfm_1 = ln_if_117_acc_itm_13_1 & (~ ln_if_118_acc_itm_14_1);
  assign ln_land_119_lpi_1_dfm_1 = ln_if_118_acc_itm_14_1 & (~ ln_if_119_acc_itm_9_1);
  assign ln_land_120_lpi_1_dfm_1 = ln_if_119_acc_itm_9_1 & (~ ln_if_120_acc_itm_14_1);
  assign ln_land_121_lpi_1_dfm_1 = ln_if_120_acc_itm_14_1 & (~ ln_if_121_acc_itm_13_1);
  assign ln_land_122_lpi_1_dfm_1 = ln_if_121_acc_itm_13_1 & (~ ln_if_122_acc_itm_14_1);
  assign ln_land_123_lpi_1_dfm_1 = ln_if_122_acc_itm_14_1 & (~ ln_if_123_acc_itm_12_1);
  assign ln_land_124_lpi_1_dfm_1 = ln_if_123_acc_itm_12_1 & (~ ln_if_124_acc_itm_14_1);
  assign ln_land_125_lpi_1_dfm_1 = ln_if_124_acc_itm_14_1 & (~ ln_if_125_acc_itm_13_1);
  assign ln_land_126_lpi_1_dfm_1 = ln_if_125_acc_itm_13_1 & (~ ln_if_126_acc_itm_14_1);
  assign ln_land_127_lpi_1_dfm_1 = ln_if_126_acc_itm_14_1 & (~ ln_if_127_acc_itm_11_1);
  assign ln_land_128_lpi_1_dfm_1 = ln_if_127_acc_itm_11_1 & (~ ln_if_128_acc_itm_14_1);
  assign ln_land_129_lpi_1_dfm_1 = ln_if_128_acc_itm_14_1 & (~ ln_if_129_acc_itm_13_1);
  assign ln_land_130_lpi_1_dfm_1 = ln_if_129_acc_itm_13_1 & (~ ln_if_130_acc_itm_14_1);
  assign ln_land_131_lpi_1_dfm_1 = ln_if_130_acc_itm_14_1 & (~ ln_if_131_acc_itm_12_1);
  assign ln_land_132_lpi_1_dfm_1 = ln_if_131_acc_itm_12_1 & (~ ln_if_132_acc_itm_14_1);
  assign ln_land_133_lpi_1_dfm_1 = ln_if_132_acc_itm_14_1 & (~ ln_if_133_acc_itm_13_1);
  assign ln_land_134_lpi_1_dfm_1 = ln_if_133_acc_itm_13_1 & (~ ln_if_134_acc_itm_14_1);
  assign ln_land_135_lpi_1_dfm_1 = ln_if_134_acc_itm_14_1 & (~ ln_if_135_acc_itm_10_1);
  assign ln_land_136_lpi_1_dfm_1 = ln_if_135_acc_itm_10_1 & (~ ln_if_136_acc_itm_14_1);
  assign ln_land_137_lpi_1_dfm_1 = ln_if_136_acc_itm_14_1 & (~ ln_if_137_acc_itm_13_1);
  assign ln_land_138_lpi_1_dfm_1 = ln_if_137_acc_itm_13_1 & (~ ln_if_138_acc_itm_14_1);
  assign ln_land_139_lpi_1_dfm_1 = ln_if_138_acc_itm_14_1 & (~ ln_if_139_acc_itm_12_1);
  assign ln_land_140_lpi_1_dfm_1 = ln_if_139_acc_itm_12_1 & (~ ln_if_140_acc_itm_14_1);
  assign ln_and_48_ssc_1 = ln_if_52_acc_itm_14_1 & (~ ln_if_53_acc_itm_14_1) & (~(ln_land_55_lpi_1_dfm_1
      | ln_land_56_lpi_1_dfm_1)) & (~(ln_land_57_lpi_1_dfm_1 | ln_land_58_lpi_1_dfm_1))
      & (~(ln_land_59_lpi_1_dfm_1 | ln_land_60_lpi_1_dfm_1)) & (~(ln_land_61_lpi_1_dfm_1
      | ln_land_62_lpi_1_dfm_1)) & (~(ln_land_63_lpi_1_dfm_1 | ln_land_64_lpi_1_dfm_1))
      & (~(ln_land_65_lpi_1_dfm_1 | ln_land_66_lpi_1_dfm_1)) & (~(ln_land_67_lpi_1_dfm_1
      | ln_land_68_lpi_1_dfm_1)) & (~(ln_land_69_lpi_1_dfm_1 | ln_land_70_lpi_1_dfm_1))
      & (~(ln_land_71_lpi_1_dfm_1 | ln_land_72_lpi_1_dfm_1)) & (~(ln_land_73_lpi_1_dfm_1
      | ln_land_74_lpi_1_dfm_1)) & (~(ln_land_75_lpi_1_dfm_1 | ln_land_76_lpi_1_dfm_1))
      & (~(ln_land_77_lpi_1_dfm_1 | ln_land_78_lpi_1_dfm_1)) & (~(ln_land_79_lpi_1_dfm_1
      | ln_land_80_lpi_1_dfm_1)) & (~(ln_land_81_lpi_1_dfm_1 | ln_land_82_lpi_1_dfm_1))
      & (~(ln_land_83_lpi_1_dfm_1 | ln_land_84_lpi_1_dfm_1)) & (~(ln_land_85_lpi_1_dfm_1
      | ln_land_86_lpi_1_dfm_1)) & (~(ln_land_87_lpi_1_dfm_1 | ln_land_88_lpi_1_dfm_1))
      & (~(ln_land_89_lpi_1_dfm_1 | ln_land_90_lpi_1_dfm_1)) & (~(ln_land_91_lpi_1_dfm_1
      | ln_land_92_lpi_1_dfm_1)) & (~(ln_land_93_lpi_1_dfm_1 | ln_land_94_lpi_1_dfm_1))
      & (~(ln_land_95_lpi_1_dfm_1 | ln_land_96_lpi_1_dfm_1)) & (~(ln_land_97_lpi_1_dfm_1
      | ln_land_98_lpi_1_dfm_1)) & (~(ln_land_99_lpi_1_dfm_1 | ln_land_100_lpi_1_dfm_1))
      & (~(ln_land_101_lpi_1_dfm_1 | ln_land_102_lpi_1_dfm_1)) & (~(ln_land_103_lpi_1_dfm_1
      | ln_land_104_lpi_1_dfm_1)) & (~(ln_land_105_lpi_1_dfm_1 | ln_land_106_lpi_1_dfm_1))
      & (~(ln_land_107_lpi_1_dfm_1 | ln_land_108_lpi_1_dfm_1)) & (~(ln_land_109_lpi_1_dfm_1
      | ln_land_110_lpi_1_dfm_1)) & (~(ln_land_111_lpi_1_dfm_1 | ln_land_112_lpi_1_dfm_1))
      & (~(ln_land_113_lpi_1_dfm_1 | ln_land_114_lpi_1_dfm_1)) & (~(ln_land_115_lpi_1_dfm_1
      | ln_land_116_lpi_1_dfm_1)) & (~(ln_land_117_lpi_1_dfm_1 | ln_land_118_lpi_1_dfm_1))
      & (~(ln_land_119_lpi_1_dfm_1 | ln_land_120_lpi_1_dfm_1)) & (~(ln_land_121_lpi_1_dfm_1
      | ln_land_122_lpi_1_dfm_1)) & (~(ln_land_123_lpi_1_dfm_1 | ln_land_124_lpi_1_dfm_1))
      & (~(ln_land_125_lpi_1_dfm_1 | ln_land_126_lpi_1_dfm_1)) & (~(ln_land_127_lpi_1_dfm_1
      | ln_land_128_lpi_1_dfm_1)) & (~(ln_land_129_lpi_1_dfm_1 | ln_land_130_lpi_1_dfm_1))
      & (~(ln_land_131_lpi_1_dfm_1 | ln_land_132_lpi_1_dfm_1)) & (~(ln_land_133_lpi_1_dfm_1
      | ln_land_134_lpi_1_dfm_1)) & (~(ln_land_135_lpi_1_dfm_1 | ln_land_136_lpi_1_dfm_1))
      & (~(ln_land_137_lpi_1_dfm_1 | ln_land_138_lpi_1_dfm_1)) & (~(ln_land_139_lpi_1_dfm_1
      | ln_land_140_lpi_1_dfm_1));
  assign ln_land_54_lpi_1_dfm_1 = ln_if_53_acc_itm_14_1 & (~ ln_if_54_acc_itm_12_1);
  assign ln_land_55_lpi_1_dfm_1 = ln_if_54_acc_itm_12_1 & (~ ln_if_55_acc_itm_14_1);
  assign ln_land_56_lpi_1_dfm_1 = ln_if_55_acc_itm_14_1 & (~ ln_if_56_acc_itm_13_1);
  assign ln_land_57_lpi_1_dfm_1 = ln_if_56_acc_itm_13_1 & (~ ln_if_57_acc_itm_14_1);
  assign ln_land_58_lpi_1_dfm_1 = ln_if_57_acc_itm_14_1 & (~ ln_if_58_acc_itm_9_1);
  assign ln_land_59_lpi_1_dfm_1 = ln_if_58_acc_itm_9_1 & (~ ln_if_59_acc_itm_14_1);
  assign ln_land_60_lpi_1_dfm_1 = ln_if_59_acc_itm_14_1 & (~ ln_if_60_acc_itm_14_1);
  assign ln_land_61_lpi_1_dfm_1 = ln_if_60_acc_itm_14_1 & (~ ln_if_61_acc_itm_13_1);
  assign ln_land_62_lpi_1_dfm_1 = ln_if_61_acc_itm_13_1 & (~ ln_if_62_acc_itm_14_1);
  assign ln_land_63_lpi_1_dfm_1 = ln_if_62_acc_itm_14_1 & (~ ln_if_63_acc_itm_10_1);
  assign ln_land_64_lpi_1_dfm_1 = ln_if_63_acc_itm_10_1 & (~ ln_if_64_acc_itm_14_1);
  assign ln_land_65_lpi_1_dfm_1 = ln_if_64_acc_itm_14_1 & (~ ln_if_65_acc_itm_13_1);
  assign ln_land_66_lpi_1_dfm_1 = ln_if_65_acc_itm_13_1 & (~ ln_if_66_acc_itm_14_1);
  assign ln_land_67_lpi_1_dfm_1 = ln_if_66_acc_itm_14_1 & (~ ln_if_67_acc_itm_14_1);
  assign ln_land_68_lpi_1_dfm_1 = ln_if_67_acc_itm_14_1 & (~ ln_if_68_acc_itm_8_1);
  assign ln_land_69_lpi_1_dfm_1 = ln_if_68_acc_itm_8_1 & (~ ln_if_69_acc_itm_14_1);
  assign ln_land_70_lpi_1_dfm_1 = ln_if_69_acc_itm_14_1 & (~ ln_if_70_acc_itm_13_1);
  assign ln_land_71_lpi_1_dfm_1 = ln_if_70_acc_itm_13_1 & (~ ln_if_71_acc_itm_14_1);
  assign ln_land_72_lpi_1_dfm_1 = ln_if_71_acc_itm_14_1 & (~ ln_if_72_acc_itm_12_1);
  assign ln_land_73_lpi_1_dfm_1 = ln_if_72_acc_itm_12_1 & (~ ln_if_73_acc_itm_14_1);
  assign ln_land_74_lpi_1_dfm_1 = ln_if_73_acc_itm_14_1 & (~ ln_if_74_acc_itm_14_1);
  assign ln_land_75_lpi_1_dfm_1 = ln_if_74_acc_itm_14_1 & (~ ln_if_75_acc_itm_13_1);
  assign ln_land_76_lpi_1_dfm_1 = ln_if_75_acc_itm_13_1 & (~ ln_if_76_acc_itm_14_1);
  assign ln_land_98_lpi_1_dfm_1 = ln_if_97_acc_itm_14_1 & (~ ln_if_98_acc_itm_13_1);
  assign ln_land_99_lpi_1_dfm_1 = ln_if_98_acc_itm_13_1 & (~ ln_if_99_acc_itm_14_1);
  assign ln_land_100_lpi_1_dfm_1 = ln_if_99_acc_itm_14_1 & (~ ln_if_100_acc_itm_12_1);
  assign ln_land_101_lpi_1_dfm_1 = ln_if_100_acc_itm_12_1 & (~ ln_if_101_acc_itm_14_1);
  assign ln_land_102_lpi_1_dfm_1 = ln_if_101_acc_itm_14_1 & (~ ln_if_102_acc_itm_14_1);
  assign ln_land_103_lpi_1_dfm_1 = ln_if_102_acc_itm_14_1 & (~ ln_if_103_acc_itm_13_1);
  assign ln_land_104_lpi_1_dfm_1 = ln_if_103_acc_itm_13_1 & (~ ln_if_104_acc_itm_14_1);
  assign ln_land_105_lpi_1_dfm_1 = ln_if_104_acc_itm_14_1 & (~ ln_if_105_acc_itm_12_1);
  assign ln_land_106_lpi_1_dfm_1 = ln_if_105_acc_itm_12_1 & (~ ln_if_106_acc_itm_14_1);
  assign ln_land_107_lpi_1_dfm_1 = ln_if_106_acc_itm_14_1 & (~ ln_if_107_acc_itm_13_1);
  assign ln_land_108_lpi_1_dfm_1 = ln_if_107_acc_itm_13_1 & (~ ln_if_108_acc_itm_14_1);
  assign ln_land_109_lpi_1_dfm_1 = ln_if_108_acc_itm_14_1 & (~ ln_if_109_acc_itm_14_1);
  assign ln_land_110_lpi_1_dfm_1 = ln_if_109_acc_itm_14_1 & (~ ln_if_110_acc_itm_12_1);
  assign ln_land_111_lpi_1_dfm_1 = ln_if_110_acc_itm_12_1 & (~ ln_if_111_acc_itm_14_1);
  assign ln_land_112_lpi_1_dfm_1 = ln_if_111_acc_itm_14_1 & (~ ln_if_112_acc_itm_13_1);
  assign ln_land_113_lpi_1_dfm_1 = ln_if_112_acc_itm_13_1 & (~ ln_if_113_acc_itm_14_1);
  assign ln_land_141_lpi_1_dfm_1 = ln_if_140_acc_itm_14_1 & (~ ln_if_141_acc_itm_13_1);
  assign ln_land_142_lpi_1_dfm_1 = ln_if_141_acc_itm_13_1 & (~ ln_if_142_acc_itm_14_1);
  assign ln_and_138_ssc_1 = ln_if_142_acc_itm_14_1 & (~ ln_if_143_acc_itm_11_1);
  assign ln_land_144_lpi_1_dfm_1 = ln_if_143_acc_itm_11_1 & (~ ln_if_144_acc_itm_14_1);
  assign ln_land_172_lpi_1_dfm_1 = ln_if_171_acc_itm_12_1 & (~ ln_if_172_acc_itm_14_1);
  assign ln_land_173_lpi_1_dfm_1 = ln_if_172_acc_itm_14_1 & (~ ln_if_173_acc_itm_13_1);
  assign ln_land_174_lpi_1_dfm_1 = ln_if_173_acc_itm_13_1 & (~ ln_if_174_acc_itm_14_1);
  assign ln_land_175_lpi_1_dfm_1 = ln_if_174_acc_itm_14_1 & (~ ln_if_175_acc_itm_11_1);
  assign ln_land_176_lpi_1_dfm_1 = ln_if_175_acc_itm_11_1 & (~ ln_if_176_acc_itm_14_1);
  assign ln_land_177_lpi_1_dfm_1 = ln_if_176_acc_itm_14_1 & (~ ln_if_177_acc_itm_13_1);
  assign ln_land_178_lpi_1_dfm_1 = ln_if_177_acc_itm_13_1 & (~ ln_if_178_acc_itm_14_1);
  assign ln_land_179_lpi_1_dfm_1 = ln_if_178_acc_itm_14_1 & (~ ln_if_179_acc_itm_12_1);
  assign ln_land_180_lpi_1_dfm_1 = ln_if_179_acc_itm_12_1 & (~ ln_if_180_acc_itm_14_1);
  assign ln_land_181_lpi_1_dfm_1 = ln_if_180_acc_itm_14_1 & (~ ln_if_181_acc_itm_13_1);
  assign ln_land_182_lpi_1_dfm_1 = ln_if_181_acc_itm_13_1 & (~ ln_if_182_acc_itm_14_1);
  assign ln_land_183_lpi_1_dfm_1 = ln_if_182_acc_itm_14_1 & (~ ln_if_183_acc_itm_9_1);
  assign ln_land_184_lpi_1_dfm_1 = ln_if_183_acc_itm_9_1 & (~ ln_if_184_acc_itm_14_1);
  assign ln_land_185_lpi_1_dfm_1 = ln_if_184_acc_itm_14_1 & (~ ln_if_185_acc_itm_13_1);
  assign ln_land_186_lpi_1_dfm_1 = ln_if_185_acc_itm_13_1 & (~ ln_if_186_acc_itm_14_1);
  assign ln_land_187_lpi_1_dfm_1 = ln_if_186_acc_itm_14_1 & (~ ln_if_187_acc_itm_12_1);
  assign ln_land_188_lpi_1_dfm_1 = ln_if_187_acc_itm_12_1 & (~ ln_if_188_acc_itm_14_1);
  assign ln_land_189_lpi_1_dfm_1 = ln_if_188_acc_itm_14_1 & (~ ln_if_189_acc_itm_13_1);
  assign ln_land_190_lpi_1_dfm_1 = ln_if_189_acc_itm_13_1 & (~ ln_if_190_acc_itm_14_1);
  assign ln_land_191_lpi_1_dfm_1 = ln_if_190_acc_itm_14_1 & (~ ln_if_191_acc_itm_11_1);
  assign ln_land_192_lpi_1_dfm_1 = ln_if_191_acc_itm_11_1 & (~ ln_if_192_acc_itm_14_1);
  assign ln_land_193_lpi_1_dfm_1 = ln_if_192_acc_itm_14_1 & (~ ln_if_193_acc_itm_13_1);
  assign ln_land_194_lpi_1_dfm_1 = ln_if_193_acc_itm_13_1 & (~ ln_if_194_acc_itm_14_1);
  assign ln_land_214_lpi_1_dfm_1 = ln_if_213_acc_itm_13_1 & (~ ln_if_214_acc_itm_14_1);
  assign ln_land_215_lpi_1_dfm_1 = ln_if_214_acc_itm_14_1 & (~ ln_if_215_acc_itm_8_1);
  assign ln_land_216_lpi_1_dfm_1 = ln_if_215_acc_itm_8_1 & (~ ln_if_216_acc_itm_14_1);
  assign ln_land_217_lpi_1_dfm_1 = ln_if_216_acc_itm_14_1 & (~ ln_if_217_acc_itm_13_1);
  assign ln_land_218_lpi_1_dfm_1 = ln_if_217_acc_itm_13_1 & (~ ln_if_218_acc_itm_14_1);
  assign ln_land_219_lpi_1_dfm_1 = ln_if_218_acc_itm_14_1 & (~ ln_if_219_acc_itm_12_1);
  assign ln_land_220_lpi_1_dfm_1 = ln_if_219_acc_itm_12_1 & (~ ln_if_220_acc_itm_14_1);
  assign ln_land_221_lpi_1_dfm_1 = ln_if_220_acc_itm_14_1 & (~ ln_if_221_acc_itm_13_1);
  assign ln_land_222_lpi_1_dfm_1 = ln_if_221_acc_itm_13_1 & (~ ln_if_222_acc_itm_14_1);
  assign ln_land_223_lpi_1_dfm_1 = ln_if_222_acc_itm_14_1 & (~ ln_if_223_acc_itm_11_1);
  assign ln_land_224_lpi_1_dfm_1 = ln_if_223_acc_itm_11_1 & (~ ln_if_224_acc_itm_14_1);
  assign ln_land_225_lpi_1_dfm_1 = ln_if_224_acc_itm_14_1 & (~ ln_if_225_acc_itm_13_1);
  assign ln_land_226_lpi_1_dfm_1 = ln_if_225_acc_itm_13_1 & (~ ln_if_226_acc_itm_14_1);
  assign ln_land_227_lpi_1_dfm_1 = ln_if_226_acc_itm_14_1 & (~ ln_if_227_acc_itm_12_1);
  assign ln_land_228_lpi_1_dfm_1 = ln_if_227_acc_itm_12_1 & (~ ln_if_228_acc_itm_14_1);
  assign ln_land_240_lpi_1_dfm_1 = ln_if_239_acc_itm_11_1 & (~ ln_if_240_acc_itm_14_1);
  assign ln_land_241_lpi_1_dfm_1 = ln_if_240_acc_itm_14_1 & (~ ln_if_241_acc_itm_13_1);
  assign ln_land_242_lpi_1_dfm_1 = ln_if_241_acc_itm_13_1 & (~ ln_if_242_acc_itm_14_1);
  assign ln_land_243_lpi_1_dfm_1 = ln_if_242_acc_itm_14_1 & (~ ln_if_243_acc_itm_12_1);
  assign ln_land_244_lpi_1_dfm_1 = ln_if_243_acc_itm_12_1 & (~ ln_if_244_acc_itm_14_1);
  assign ln_and_140_ssc_1 = ln_if_144_acc_itm_14_1 & (~ ln_if_145_acc_itm_13_1) &
      (~(ln_land_147_lpi_1_dfm_1 | ln_land_148_lpi_1_dfm_1)) & (~(ln_land_149_lpi_1_dfm_1
      | ln_land_150_lpi_1_dfm_1)) & (~(ln_land_151_lpi_1_dfm_1 | ln_land_152_lpi_1_dfm_1))
      & (~(ln_land_153_lpi_1_dfm_1 | ln_land_154_lpi_1_dfm_1)) & (~(ln_land_155_lpi_1_dfm_1
      | ln_land_156_lpi_1_dfm_1)) & (~(ln_land_157_lpi_1_dfm_1 | ln_land_158_lpi_1_dfm_1))
      & (~(ln_land_159_lpi_1_dfm_1 | ln_land_160_lpi_1_dfm_1)) & (~(ln_land_161_lpi_1_dfm_1
      | ln_land_162_lpi_1_dfm_1)) & (~(ln_land_163_lpi_1_dfm_1 | ln_land_164_lpi_1_dfm_1))
      & (~(ln_land_165_lpi_1_dfm_1 | ln_land_166_lpi_1_dfm_1)) & (~(ln_land_167_lpi_1_dfm_1
      | ln_land_168_lpi_1_dfm_1)) & (~(ln_land_169_lpi_1_dfm_1 | ln_land_170_lpi_1_dfm_1))
      & (~(ln_land_171_lpi_1_dfm_1 | ln_land_172_lpi_1_dfm_1)) & (~(ln_land_173_lpi_1_dfm_1
      | ln_land_174_lpi_1_dfm_1)) & (~(ln_land_175_lpi_1_dfm_1 | ln_land_176_lpi_1_dfm_1))
      & (~(ln_land_177_lpi_1_dfm_1 | ln_land_178_lpi_1_dfm_1)) & (~(ln_land_179_lpi_1_dfm_1
      | ln_land_180_lpi_1_dfm_1)) & (~(ln_land_181_lpi_1_dfm_1 | ln_land_182_lpi_1_dfm_1))
      & (~(ln_land_183_lpi_1_dfm_1 | ln_land_184_lpi_1_dfm_1)) & (~(ln_land_185_lpi_1_dfm_1
      | ln_land_186_lpi_1_dfm_1)) & (~(ln_land_187_lpi_1_dfm_1 | ln_land_188_lpi_1_dfm_1))
      & (~(ln_land_189_lpi_1_dfm_1 | ln_land_190_lpi_1_dfm_1)) & (~(ln_land_191_lpi_1_dfm_1
      | ln_land_192_lpi_1_dfm_1)) & (~(ln_land_193_lpi_1_dfm_1 | ln_land_194_lpi_1_dfm_1))
      & (~(ln_land_195_lpi_1_dfm_1 | ln_land_196_lpi_1_dfm_1)) & (~(ln_land_197_lpi_1_dfm_1
      | ln_land_198_lpi_1_dfm_1)) & (~(ln_land_199_lpi_1_dfm_1 | ln_land_200_lpi_1_dfm_1))
      & (~(ln_land_201_lpi_1_dfm_1 | ln_land_202_lpi_1_dfm_1)) & (~(ln_land_203_lpi_1_dfm_1
      | ln_land_204_lpi_1_dfm_1)) & (~(ln_land_205_lpi_1_dfm_1 | ln_land_206_lpi_1_dfm_1))
      & (~(ln_land_207_lpi_1_dfm_1 | ln_land_208_lpi_1_dfm_1)) & (~(ln_land_209_lpi_1_dfm_1
      | ln_land_210_lpi_1_dfm_1)) & (~(ln_land_211_lpi_1_dfm_1 | ln_land_212_lpi_1_dfm_1))
      & (~(ln_land_213_lpi_1_dfm_1 | ln_land_214_lpi_1_dfm_1)) & (~(ln_land_215_lpi_1_dfm_1
      | ln_land_216_lpi_1_dfm_1)) & (~(ln_land_217_lpi_1_dfm_1 | ln_land_218_lpi_1_dfm_1))
      & (~(ln_land_219_lpi_1_dfm_1 | ln_land_220_lpi_1_dfm_1)) & (~(ln_land_221_lpi_1_dfm_1
      | ln_land_222_lpi_1_dfm_1)) & (~(ln_land_223_lpi_1_dfm_1 | ln_land_224_lpi_1_dfm_1))
      & (~(ln_land_225_lpi_1_dfm_1 | ln_land_226_lpi_1_dfm_1)) & (~(ln_land_227_lpi_1_dfm_1
      | ln_land_228_lpi_1_dfm_1)) & ln_and_368_m1c_1;
  assign ln_land_146_lpi_1_dfm_1 = ln_if_145_acc_itm_13_1 & (~ ln_if_146_acc_itm_14_1);
  assign ln_land_147_lpi_1_dfm_1 = ln_if_146_acc_itm_14_1 & (~ ln_if_147_acc_itm_12_1);
  assign ln_land_148_lpi_1_dfm_1 = ln_if_147_acc_itm_12_1 & (~ ln_if_148_acc_itm_14_1);
  assign ln_land_149_lpi_1_dfm_1 = ln_if_148_acc_itm_14_1 & (~ ln_if_149_acc_itm_13_1);
  assign ln_land_150_lpi_1_dfm_1 = ln_if_149_acc_itm_13_1 & (~ ln_if_150_acc_itm_14_1);
  assign ln_land_151_lpi_1_dfm_1 = ln_if_150_acc_itm_14_1 & (~ ln_if_151_acc_itm_7_1);
  assign ln_land_152_lpi_1_dfm_1 = ln_if_151_acc_itm_7_1 & (~ ln_if_152_acc_itm_14_1);
  assign ln_land_153_lpi_1_dfm_1 = ln_if_152_acc_itm_14_1 & (~ ln_if_153_acc_itm_13_1);
  assign ln_land_154_lpi_1_dfm_1 = ln_if_153_acc_itm_13_1 & (~ ln_if_154_acc_itm_14_1);
  assign ln_land_155_lpi_1_dfm_1 = ln_if_154_acc_itm_14_1 & (~ ln_if_155_acc_itm_12_1);
  assign ln_land_156_lpi_1_dfm_1 = ln_if_155_acc_itm_12_1 & (~ ln_if_156_acc_itm_14_1);
  assign ln_land_157_lpi_1_dfm_1 = ln_if_156_acc_itm_14_1 & (~ ln_if_157_acc_itm_13_1);
  assign ln_land_158_lpi_1_dfm_1 = ln_if_157_acc_itm_13_1 & (~ ln_if_158_acc_itm_14_1);
  assign ln_land_159_lpi_1_dfm_1 = ln_if_158_acc_itm_14_1 & (~ ln_if_159_acc_itm_11_1);
  assign ln_land_160_lpi_1_dfm_1 = ln_if_159_acc_itm_11_1 & (~ ln_if_160_acc_itm_14_1);
  assign ln_land_161_lpi_1_dfm_1 = ln_if_160_acc_itm_14_1 & (~ ln_if_161_acc_itm_13_1);
  assign ln_land_162_lpi_1_dfm_1 = ln_if_161_acc_itm_13_1 & (~ ln_if_162_acc_itm_14_1);
  assign ln_land_163_lpi_1_dfm_1 = ln_if_162_acc_itm_14_1 & (~ ln_if_163_acc_itm_12_1);
  assign ln_land_164_lpi_1_dfm_1 = ln_if_163_acc_itm_12_1 & (~ ln_if_164_acc_itm_14_1);
  assign ln_land_165_lpi_1_dfm_1 = ln_if_164_acc_itm_14_1 & (~ ln_if_165_acc_itm_13_1);
  assign ln_land_166_lpi_1_dfm_1 = ln_if_165_acc_itm_13_1 & (~ ln_if_166_acc_itm_14_1);
  assign ln_land_167_lpi_1_dfm_1 = ln_if_166_acc_itm_14_1 & (~ ln_if_167_acc_itm_10_1);
  assign ln_land_168_lpi_1_dfm_1 = ln_if_167_acc_itm_10_1 & (~ ln_if_168_acc_itm_14_1);
  assign ln_land_169_lpi_1_dfm_1 = ln_if_168_acc_itm_14_1 & (~ ln_if_169_acc_itm_13_1);
  assign ln_land_170_lpi_1_dfm_1 = ln_if_169_acc_itm_13_1 & (~ ln_if_170_acc_itm_14_1);
  assign ln_land_171_lpi_1_dfm_1 = ln_if_170_acc_itm_14_1 & (~ ln_if_171_acc_itm_12_1);
  assign ln_land_195_lpi_1_dfm_1 = ln_if_194_acc_itm_14_1 & (~ ln_if_195_acc_itm_12_1);
  assign ln_land_196_lpi_1_dfm_1 = ln_if_195_acc_itm_12_1 & (~ ln_if_196_acc_itm_14_1);
  assign ln_land_197_lpi_1_dfm_1 = ln_if_196_acc_itm_14_1 & (~ ln_if_197_acc_itm_13_1);
  assign ln_land_198_lpi_1_dfm_1 = ln_if_197_acc_itm_13_1 & (~ ln_if_198_acc_itm_14_1);
  assign ln_land_199_lpi_1_dfm_1 = ln_if_198_acc_itm_14_1 & (~ ln_if_199_acc_itm_10_1);
  assign ln_land_200_lpi_1_dfm_1 = ln_if_199_acc_itm_10_1 & (~ ln_if_200_acc_itm_14_1);
  assign ln_land_201_lpi_1_dfm_1 = ln_if_200_acc_itm_14_1 & (~ ln_if_201_acc_itm_13_1);
  assign ln_land_202_lpi_1_dfm_1 = ln_if_201_acc_itm_13_1 & (~ ln_if_202_acc_itm_14_1);
  assign ln_land_203_lpi_1_dfm_1 = ln_if_202_acc_itm_14_1 & (~ ln_if_203_acc_itm_12_1);
  assign ln_land_204_lpi_1_dfm_1 = ln_if_203_acc_itm_12_1 & (~ ln_if_204_acc_itm_14_1);
  assign ln_land_205_lpi_1_dfm_1 = ln_if_204_acc_itm_14_1 & (~ ln_if_205_acc_itm_13_1);
  assign ln_land_206_lpi_1_dfm_1 = ln_if_205_acc_itm_13_1 & (~ ln_if_206_acc_itm_14_1);
  assign ln_land_207_lpi_1_dfm_1 = ln_if_206_acc_itm_14_1 & (~ ln_if_207_acc_itm_11_1);
  assign ln_land_208_lpi_1_dfm_1 = ln_if_207_acc_itm_11_1 & (~ ln_if_208_acc_itm_14_1);
  assign ln_land_209_lpi_1_dfm_1 = ln_if_208_acc_itm_14_1 & (~ ln_if_209_acc_itm_13_1);
  assign ln_land_210_lpi_1_dfm_1 = ln_if_209_acc_itm_13_1 & (~ ln_if_210_acc_itm_14_1);
  assign ln_land_211_lpi_1_dfm_1 = ln_if_210_acc_itm_14_1 & (~ ln_if_211_acc_itm_12_1);
  assign ln_land_212_lpi_1_dfm_1 = ln_if_211_acc_itm_12_1 & (~ ln_if_212_acc_itm_14_1);
  assign ln_land_213_lpi_1_dfm_1 = ln_if_212_acc_itm_14_1 & (~ ln_if_213_acc_itm_13_1);
  assign ln_land_229_lpi_1_dfm_1 = ln_if_228_acc_itm_14_1 & (~ ln_if_229_acc_itm_13_1);
  assign ln_land_230_lpi_1_dfm_1 = ln_if_229_acc_itm_13_1 & (~ ln_if_230_acc_itm_14_1);
  assign ln_land_231_lpi_1_dfm_1 = ln_if_230_acc_itm_14_1 & (~ ln_if_231_acc_itm_10_1);
  assign ln_land_232_lpi_1_dfm_1 = ln_if_231_acc_itm_10_1 & (~ ln_if_232_acc_itm_14_1);
  assign ln_land_233_lpi_1_dfm_1 = ln_if_232_acc_itm_14_1 & (~ ln_if_233_acc_itm_13_1);
  assign ln_land_234_lpi_1_dfm_1 = ln_if_233_acc_itm_13_1 & (~ ln_if_234_acc_itm_14_1);
  assign ln_land_235_lpi_1_dfm_1 = ln_if_234_acc_itm_14_1 & (~ ln_if_235_acc_itm_12_1);
  assign ln_land_236_lpi_1_dfm_1 = ln_if_235_acc_itm_12_1 & (~ ln_if_236_acc_itm_14_1);
  assign ln_land_237_lpi_1_dfm_1 = ln_if_236_acc_itm_14_1 & (~ ln_if_237_acc_itm_13_1);
  assign ln_land_238_lpi_1_dfm_1 = ln_if_237_acc_itm_13_1 & (~ ln_if_238_acc_itm_14_1);
  assign ln_land_239_lpi_1_dfm_1 = ln_if_238_acc_itm_14_1 & (~ ln_if_239_acc_itm_11_1);
  assign nl_ln_if_252_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111111101;
  assign ln_if_252_acc_nl = nl_ln_if_252_acc_nl[12:0];
  assign ln_if_252_acc_itm_12_1 = readslicef_13_1_12(ln_if_252_acc_nl);
  assign nl_ln_if_244_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111111011101;
  assign ln_if_244_acc_nl = nl_ln_if_244_acc_nl[14:0];
  assign ln_if_244_acc_itm_14_1 = readslicef_15_1_14(ln_if_244_acc_nl);
  assign nl_ln_if_245_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111101111;
  assign ln_if_245_acc_nl = nl_ln_if_245_acc_nl[13:0];
  assign ln_if_245_acc_itm_13_1 = readslicef_14_1_13(ln_if_245_acc_nl);
  assign nl_ln_if_251_acc_nl = conv_u2u_10_11(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:4])
      + 11'b11111111111;
  assign ln_if_251_acc_nl = nl_ln_if_251_acc_nl[10:0];
  assign ln_if_251_acc_itm_10_1 = readslicef_11_1_10(ln_if_251_acc_nl);
  assign nl_ln_if_250_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111111011;
  assign ln_if_250_acc_nl = nl_ln_if_250_acc_nl[12:0];
  assign ln_if_250_acc_itm_12_1 = readslicef_13_1_12(ln_if_250_acc_nl);
  assign nl_ln_if_249_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:3])
      + 12'b111111111101;
  assign ln_if_249_acc_nl = nl_ln_if_249_acc_nl[11:0];
  assign ln_if_249_acc_itm_11_1 = readslicef_12_1_11(ln_if_249_acc_nl);
  assign nl_ln_if_248_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111111001;
  assign ln_if_248_acc_nl = nl_ln_if_248_acc_nl[12:0];
  assign ln_if_248_acc_itm_12_1 = readslicef_13_1_12(ln_if_248_acc_nl);
  assign nl_ln_if_247_acc_nl = conv_u2u_9_10(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:5])
      + 10'b1111111111;
  assign ln_if_247_acc_nl = nl_ln_if_247_acc_nl[9:0];
  assign ln_if_247_acc_itm_9_1 = readslicef_10_1_9(ln_if_247_acc_nl);
  assign nl_ln_if_246_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111111011111;
  assign ln_if_246_acc_nl = nl_ln_if_246_acc_nl[14:0];
  assign ln_if_246_acc_itm_14_1 = readslicef_15_1_14(ln_if_246_acc_nl);
  assign ln_nor_3_cse_1 = ~(ln_and_138_ssc_1 | ln_land_144_lpi_1_dfm_1);
  assign ln_nor_1_cse_1 = ~(ln_and_2_ssc_1 | ln_land_6_lpi_1_dfm_1);
  assign ln_land_8_lpi_1_dfm_1 = ln_if_7_acc_itm_5_1 & (~ ln_if_8_acc_itm_14_1);
  assign ln_land_9_lpi_1_dfm_1 = ln_if_8_acc_itm_14_1 & (~ ln_if_9_acc_itm_13_1);
  assign ln_land_11_lpi_1_dfm_1 = ln_if_10_acc_itm_14_1 & (~ ln_if_11_acc_itm_14_1);
  assign ln_land_13_lpi_1_dfm_1 = ln_if_12_acc_itm_10_1 & (~ ln_if_13_acc_itm_14_1);
  assign ln_land_15_lpi_1_dfm_1 = ln_if_14_acc_itm_13_1 & (~ ln_if_15_acc_itm_14_1);
  assign ln_and_4_ssc_1 = ln_if_6_acc_itm_8_1 & (~ ln_if_7_acc_itm_5_1) & (~(ln_land_9_lpi_1_dfm_1
      | ln_land_10_lpi_1_dfm_1)) & (~(ln_land_11_lpi_1_dfm_1 | ln_land_12_lpi_1_dfm_1))
      & (~(ln_land_13_lpi_1_dfm_1 | ln_land_14_lpi_1_dfm_1)) & (~(ln_land_15_lpi_1_dfm_1
      | ln_land_16_lpi_1_dfm_1)) & (~(ln_land_17_lpi_1_dfm_1 | ln_land_18_lpi_1_dfm_1))
      & (~(ln_land_19_lpi_1_dfm_1 | ln_land_20_lpi_1_dfm_1)) & (~(ln_land_21_lpi_1_dfm_1
      | ln_land_22_lpi_1_dfm_1)) & (~(ln_land_23_lpi_1_dfm_1 | ln_land_24_lpi_1_dfm_1))
      & (~(ln_land_25_lpi_1_dfm_1 | ln_land_26_lpi_1_dfm_1)) & (~(ln_land_27_lpi_1_dfm_1
      | ln_land_28_lpi_1_dfm_1)) & (~(ln_land_29_lpi_1_dfm_1 | ln_land_30_lpi_1_dfm_1))
      & (~(ln_land_31_lpi_1_dfm_1 | ln_land_32_lpi_1_dfm_1)) & (~(ln_land_33_lpi_1_dfm_1
      | ln_land_34_lpi_1_dfm_1)) & (~(ln_land_35_lpi_1_dfm_1 | ln_land_36_lpi_1_dfm_1))
      & (~(ln_land_37_lpi_1_dfm_1 | ln_land_38_lpi_1_dfm_1)) & (~(ln_land_39_lpi_1_dfm_1
      | ln_land_40_lpi_1_dfm_1)) & (~(ln_land_41_lpi_1_dfm_1 | ln_land_42_lpi_1_dfm_1))
      & (~(ln_land_43_lpi_1_dfm_1 | ln_land_44_lpi_1_dfm_1)) & (~(ln_land_45_lpi_1_dfm_1
      | ln_land_46_lpi_1_dfm_1)) & (~(ln_land_47_lpi_1_dfm_1 | ln_land_48_lpi_1_dfm_1
      | ln_land_49_lpi_1_dfm_1));
  assign ln_land_10_lpi_1_dfm_1 = ln_if_9_acc_itm_13_1 & (~ ln_if_10_acc_itm_14_1);
  assign ln_land_12_lpi_1_dfm_1 = ln_if_11_acc_itm_14_1 & (~ ln_if_12_acc_itm_10_1);
  assign ln_land_14_lpi_1_dfm_1 = ln_if_13_acc_itm_14_1 & (~ ln_if_14_acc_itm_13_1);
  assign ln_land_16_lpi_1_dfm_1 = ln_if_15_acc_itm_14_1 & (~ ln_if_16_acc_itm_12_1);
  assign ln_and_368_m1c_1 = (~(ln_land_229_lpi_1_dfm_1 | ln_land_230_lpi_1_dfm_1))
      & (~(ln_land_231_lpi_1_dfm_1 | ln_land_232_lpi_1_dfm_1)) & (~(ln_land_233_lpi_1_dfm_1
      | ln_land_234_lpi_1_dfm_1)) & (~(ln_land_235_lpi_1_dfm_1 | ln_land_236_lpi_1_dfm_1))
      & (~(ln_land_237_lpi_1_dfm_1 | ln_land_238_lpi_1_dfm_1)) & (~(ln_land_239_lpi_1_dfm_1
      | ln_land_240_lpi_1_dfm_1)) & (~(ln_land_241_lpi_1_dfm_1 | ln_land_242_lpi_1_dfm_1))
      & (~(ln_land_243_lpi_1_dfm_1 | ln_land_244_lpi_1_dfm_1));
  assign ln_land_4_lpi_1_dfm_1 = ln_if_3_acc_itm_6_1 & (~ ln_if_4_acc_itm_8_1);
  assign ln_and_2_ssc_1 = ln_if_4_acc_itm_8_1 & (~ ln_if_5_acc_itm_7_1);
  assign ln_land_6_lpi_1_dfm_1 = ln_if_5_acc_itm_7_1 & (~ ln_if_6_acc_itm_8_1);
  assign ln_nor_5_cse_1 = ~(ln_land_3_lpi_1_dfm_1 | ln_land_4_lpi_1_dfm_1);
  assign nl_ln_if_1_acc_nl = conv_u2u_7_8(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:7])
      + 8'b11111001;
  assign ln_if_1_acc_nl = nl_ln_if_1_acc_nl[7:0];
  assign ln_ret_13_0_lpi_1_dfm_258 = (readslicef_8_1_7(ln_if_1_acc_nl)) & (~ ln_if_2_acc_itm_8_1);
  assign ln_land_3_lpi_1_dfm_1 = ln_if_2_acc_itm_8_1 & (~ ln_if_3_acc_itm_6_1);
  assign ln_ln_ln_nor_8_cse_1 = ~(ln_ret_13_0_lpi_1_dfm_258 | ln_land_4_lpi_1_dfm_1);
  assign nl_ln_if_144_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101111001;
  assign ln_if_144_acc_nl = nl_ln_if_144_acc_nl[14:0];
  assign ln_if_144_acc_itm_14_1 = readslicef_15_1_14(ln_if_144_acc_nl);
  assign nl_ln_if_145_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111110111101;
  assign ln_if_145_acc_nl = nl_ln_if_145_acc_nl[13:0];
  assign ln_if_145_acc_itm_13_1 = readslicef_14_1_13(ln_if_145_acc_nl);
  assign nl_ln_if_243_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111110111;
  assign ln_if_243_acc_nl = nl_ln_if_243_acc_nl[12:0];
  assign ln_if_243_acc_itm_12_1 = readslicef_13_1_12(ln_if_243_acc_nl);
  assign nl_ln_if_242_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111111011011;
  assign ln_if_242_acc_nl = nl_ln_if_242_acc_nl[14:0];
  assign ln_if_242_acc_itm_14_1 = readslicef_15_1_14(ln_if_242_acc_nl);
  assign nl_ln_if_241_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111101101;
  assign ln_if_241_acc_nl = nl_ln_if_241_acc_nl[13:0];
  assign ln_if_241_acc_itm_13_1 = readslicef_14_1_13(ln_if_241_acc_nl);
  assign nl_ln_if_240_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111111011001;
  assign ln_if_240_acc_nl = nl_ln_if_240_acc_nl[14:0];
  assign ln_if_240_acc_itm_14_1 = readslicef_15_1_14(ln_if_240_acc_nl);
  assign nl_ln_if_239_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:3])
      + 12'b111111111011;
  assign ln_if_239_acc_nl = nl_ln_if_239_acc_nl[11:0];
  assign ln_if_239_acc_itm_11_1 = readslicef_12_1_11(ln_if_239_acc_nl);
  assign nl_ln_if_238_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111111010111;
  assign ln_if_238_acc_nl = nl_ln_if_238_acc_nl[14:0];
  assign ln_if_238_acc_itm_14_1 = readslicef_15_1_14(ln_if_238_acc_nl);
  assign nl_ln_if_237_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111101011;
  assign ln_if_237_acc_nl = nl_ln_if_237_acc_nl[13:0];
  assign ln_if_237_acc_itm_13_1 = readslicef_14_1_13(ln_if_237_acc_nl);
  assign nl_ln_if_236_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111111010101;
  assign ln_if_236_acc_nl = nl_ln_if_236_acc_nl[14:0];
  assign ln_if_236_acc_itm_14_1 = readslicef_15_1_14(ln_if_236_acc_nl);
  assign nl_ln_if_235_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111110101;
  assign ln_if_235_acc_nl = nl_ln_if_235_acc_nl[12:0];
  assign ln_if_235_acc_itm_12_1 = readslicef_13_1_12(ln_if_235_acc_nl);
  assign nl_ln_if_234_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111111010011;
  assign ln_if_234_acc_nl = nl_ln_if_234_acc_nl[14:0];
  assign ln_if_234_acc_itm_14_1 = readslicef_15_1_14(ln_if_234_acc_nl);
  assign nl_ln_if_233_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111101001;
  assign ln_if_233_acc_nl = nl_ln_if_233_acc_nl[13:0];
  assign ln_if_233_acc_itm_13_1 = readslicef_14_1_13(ln_if_233_acc_nl);
  assign nl_ln_if_232_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111111010001;
  assign ln_if_232_acc_nl = nl_ln_if_232_acc_nl[14:0];
  assign ln_if_232_acc_itm_14_1 = readslicef_15_1_14(ln_if_232_acc_nl);
  assign nl_ln_if_231_acc_nl = conv_u2u_10_11(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:4])
      + 11'b11111111101;
  assign ln_if_231_acc_nl = nl_ln_if_231_acc_nl[10:0];
  assign ln_if_231_acc_itm_10_1 = readslicef_11_1_10(ln_if_231_acc_nl);
  assign nl_ln_if_230_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111111001111;
  assign ln_if_230_acc_nl = nl_ln_if_230_acc_nl[14:0];
  assign ln_if_230_acc_itm_14_1 = readslicef_15_1_14(ln_if_230_acc_nl);
  assign nl_ln_if_229_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111100111;
  assign ln_if_229_acc_nl = nl_ln_if_229_acc_nl[13:0];
  assign ln_if_229_acc_itm_13_1 = readslicef_14_1_13(ln_if_229_acc_nl);
  assign nl_ln_if_228_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111111001101;
  assign ln_if_228_acc_nl = nl_ln_if_228_acc_nl[14:0];
  assign ln_if_228_acc_itm_14_1 = readslicef_15_1_14(ln_if_228_acc_nl);
  assign nl_ln_if_227_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111110011;
  assign ln_if_227_acc_nl = nl_ln_if_227_acc_nl[12:0];
  assign ln_if_227_acc_itm_12_1 = readslicef_13_1_12(ln_if_227_acc_nl);
  assign nl_ln_if_226_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111111001011;
  assign ln_if_226_acc_nl = nl_ln_if_226_acc_nl[14:0];
  assign ln_if_226_acc_itm_14_1 = readslicef_15_1_14(ln_if_226_acc_nl);
  assign nl_ln_if_225_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111100101;
  assign ln_if_225_acc_nl = nl_ln_if_225_acc_nl[13:0];
  assign ln_if_225_acc_itm_13_1 = readslicef_14_1_13(ln_if_225_acc_nl);
  assign nl_ln_if_224_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111111001001;
  assign ln_if_224_acc_nl = nl_ln_if_224_acc_nl[14:0];
  assign ln_if_224_acc_itm_14_1 = readslicef_15_1_14(ln_if_224_acc_nl);
  assign nl_ln_if_223_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:3])
      + 12'b111111111001;
  assign ln_if_223_acc_nl = nl_ln_if_223_acc_nl[11:0];
  assign ln_if_223_acc_itm_11_1 = readslicef_12_1_11(ln_if_223_acc_nl);
  assign nl_ln_if_222_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111111000111;
  assign ln_if_222_acc_nl = nl_ln_if_222_acc_nl[14:0];
  assign ln_if_222_acc_itm_14_1 = readslicef_15_1_14(ln_if_222_acc_nl);
  assign nl_ln_if_221_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111100011;
  assign ln_if_221_acc_nl = nl_ln_if_221_acc_nl[13:0];
  assign ln_if_221_acc_itm_13_1 = readslicef_14_1_13(ln_if_221_acc_nl);
  assign nl_ln_if_220_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111111000101;
  assign ln_if_220_acc_nl = nl_ln_if_220_acc_nl[14:0];
  assign ln_if_220_acc_itm_14_1 = readslicef_15_1_14(ln_if_220_acc_nl);
  assign nl_ln_if_219_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111110001;
  assign ln_if_219_acc_nl = nl_ln_if_219_acc_nl[12:0];
  assign ln_if_219_acc_itm_12_1 = readslicef_13_1_12(ln_if_219_acc_nl);
  assign nl_ln_if_218_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111111000011;
  assign ln_if_218_acc_nl = nl_ln_if_218_acc_nl[14:0];
  assign ln_if_218_acc_itm_14_1 = readslicef_15_1_14(ln_if_218_acc_nl);
  assign nl_ln_if_217_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111100001;
  assign ln_if_217_acc_nl = nl_ln_if_217_acc_nl[13:0];
  assign ln_if_217_acc_itm_13_1 = readslicef_14_1_13(ln_if_217_acc_nl);
  assign nl_ln_if_216_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111111000001;
  assign ln_if_216_acc_nl = nl_ln_if_216_acc_nl[14:0];
  assign ln_if_216_acc_itm_14_1 = readslicef_15_1_14(ln_if_216_acc_nl);
  assign nl_ln_if_215_acc_nl = conv_u2u_8_9(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:6])
      + 9'b111111111;
  assign ln_if_215_acc_nl = nl_ln_if_215_acc_nl[8:0];
  assign ln_if_215_acc_itm_8_1 = readslicef_9_1_8(ln_if_215_acc_nl);
  assign nl_ln_if_214_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110111111;
  assign ln_if_214_acc_nl = nl_ln_if_214_acc_nl[14:0];
  assign ln_if_214_acc_itm_14_1 = readslicef_15_1_14(ln_if_214_acc_nl);
  assign nl_ln_if_213_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111011111;
  assign ln_if_213_acc_nl = nl_ln_if_213_acc_nl[13:0];
  assign ln_if_213_acc_itm_13_1 = readslicef_14_1_13(ln_if_213_acc_nl);
  assign nl_ln_if_212_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110111101;
  assign ln_if_212_acc_nl = nl_ln_if_212_acc_nl[14:0];
  assign ln_if_212_acc_itm_14_1 = readslicef_15_1_14(ln_if_212_acc_nl);
  assign nl_ln_if_211_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111101111;
  assign ln_if_211_acc_nl = nl_ln_if_211_acc_nl[12:0];
  assign ln_if_211_acc_itm_12_1 = readslicef_13_1_12(ln_if_211_acc_nl);
  assign nl_ln_if_210_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110111011;
  assign ln_if_210_acc_nl = nl_ln_if_210_acc_nl[14:0];
  assign ln_if_210_acc_itm_14_1 = readslicef_15_1_14(ln_if_210_acc_nl);
  assign nl_ln_if_209_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111011101;
  assign ln_if_209_acc_nl = nl_ln_if_209_acc_nl[13:0];
  assign ln_if_209_acc_itm_13_1 = readslicef_14_1_13(ln_if_209_acc_nl);
  assign nl_ln_if_208_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110111001;
  assign ln_if_208_acc_nl = nl_ln_if_208_acc_nl[14:0];
  assign ln_if_208_acc_itm_14_1 = readslicef_15_1_14(ln_if_208_acc_nl);
  assign nl_ln_if_207_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:3])
      + 12'b111111110111;
  assign ln_if_207_acc_nl = nl_ln_if_207_acc_nl[11:0];
  assign ln_if_207_acc_itm_11_1 = readslicef_12_1_11(ln_if_207_acc_nl);
  assign nl_ln_if_206_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110110111;
  assign ln_if_206_acc_nl = nl_ln_if_206_acc_nl[14:0];
  assign ln_if_206_acc_itm_14_1 = readslicef_15_1_14(ln_if_206_acc_nl);
  assign nl_ln_if_205_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111011011;
  assign ln_if_205_acc_nl = nl_ln_if_205_acc_nl[13:0];
  assign ln_if_205_acc_itm_13_1 = readslicef_14_1_13(ln_if_205_acc_nl);
  assign nl_ln_if_204_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110110101;
  assign ln_if_204_acc_nl = nl_ln_if_204_acc_nl[14:0];
  assign ln_if_204_acc_itm_14_1 = readslicef_15_1_14(ln_if_204_acc_nl);
  assign nl_ln_if_203_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111101101;
  assign ln_if_203_acc_nl = nl_ln_if_203_acc_nl[12:0];
  assign ln_if_203_acc_itm_12_1 = readslicef_13_1_12(ln_if_203_acc_nl);
  assign nl_ln_if_202_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110110011;
  assign ln_if_202_acc_nl = nl_ln_if_202_acc_nl[14:0];
  assign ln_if_202_acc_itm_14_1 = readslicef_15_1_14(ln_if_202_acc_nl);
  assign nl_ln_if_201_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111011001;
  assign ln_if_201_acc_nl = nl_ln_if_201_acc_nl[13:0];
  assign ln_if_201_acc_itm_13_1 = readslicef_14_1_13(ln_if_201_acc_nl);
  assign nl_ln_if_200_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110110001;
  assign ln_if_200_acc_nl = nl_ln_if_200_acc_nl[14:0];
  assign ln_if_200_acc_itm_14_1 = readslicef_15_1_14(ln_if_200_acc_nl);
  assign nl_ln_if_199_acc_nl = conv_u2u_10_11(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:4])
      + 11'b11111111011;
  assign ln_if_199_acc_nl = nl_ln_if_199_acc_nl[10:0];
  assign ln_if_199_acc_itm_10_1 = readslicef_11_1_10(ln_if_199_acc_nl);
  assign nl_ln_if_198_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110101111;
  assign ln_if_198_acc_nl = nl_ln_if_198_acc_nl[14:0];
  assign ln_if_198_acc_itm_14_1 = readslicef_15_1_14(ln_if_198_acc_nl);
  assign nl_ln_if_197_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111010111;
  assign ln_if_197_acc_nl = nl_ln_if_197_acc_nl[13:0];
  assign ln_if_197_acc_itm_13_1 = readslicef_14_1_13(ln_if_197_acc_nl);
  assign nl_ln_if_196_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110101101;
  assign ln_if_196_acc_nl = nl_ln_if_196_acc_nl[14:0];
  assign ln_if_196_acc_itm_14_1 = readslicef_15_1_14(ln_if_196_acc_nl);
  assign nl_ln_if_195_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111101011;
  assign ln_if_195_acc_nl = nl_ln_if_195_acc_nl[12:0];
  assign ln_if_195_acc_itm_12_1 = readslicef_13_1_12(ln_if_195_acc_nl);
  assign nl_ln_if_194_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110101011;
  assign ln_if_194_acc_nl = nl_ln_if_194_acc_nl[14:0];
  assign ln_if_194_acc_itm_14_1 = readslicef_15_1_14(ln_if_194_acc_nl);
  assign nl_ln_if_193_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111010101;
  assign ln_if_193_acc_nl = nl_ln_if_193_acc_nl[13:0];
  assign ln_if_193_acc_itm_13_1 = readslicef_14_1_13(ln_if_193_acc_nl);
  assign nl_ln_if_192_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110101001;
  assign ln_if_192_acc_nl = nl_ln_if_192_acc_nl[14:0];
  assign ln_if_192_acc_itm_14_1 = readslicef_15_1_14(ln_if_192_acc_nl);
  assign nl_ln_if_191_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:3])
      + 12'b111111110101;
  assign ln_if_191_acc_nl = nl_ln_if_191_acc_nl[11:0];
  assign ln_if_191_acc_itm_11_1 = readslicef_12_1_11(ln_if_191_acc_nl);
  assign nl_ln_if_190_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110100111;
  assign ln_if_190_acc_nl = nl_ln_if_190_acc_nl[14:0];
  assign ln_if_190_acc_itm_14_1 = readslicef_15_1_14(ln_if_190_acc_nl);
  assign nl_ln_if_189_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111010011;
  assign ln_if_189_acc_nl = nl_ln_if_189_acc_nl[13:0];
  assign ln_if_189_acc_itm_13_1 = readslicef_14_1_13(ln_if_189_acc_nl);
  assign nl_ln_if_188_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110100101;
  assign ln_if_188_acc_nl = nl_ln_if_188_acc_nl[14:0];
  assign ln_if_188_acc_itm_14_1 = readslicef_15_1_14(ln_if_188_acc_nl);
  assign nl_ln_if_187_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111101001;
  assign ln_if_187_acc_nl = nl_ln_if_187_acc_nl[12:0];
  assign ln_if_187_acc_itm_12_1 = readslicef_13_1_12(ln_if_187_acc_nl);
  assign nl_ln_if_186_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110100011;
  assign ln_if_186_acc_nl = nl_ln_if_186_acc_nl[14:0];
  assign ln_if_186_acc_itm_14_1 = readslicef_15_1_14(ln_if_186_acc_nl);
  assign nl_ln_if_185_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111010001;
  assign ln_if_185_acc_nl = nl_ln_if_185_acc_nl[13:0];
  assign ln_if_185_acc_itm_13_1 = readslicef_14_1_13(ln_if_185_acc_nl);
  assign nl_ln_if_184_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110100001;
  assign ln_if_184_acc_nl = nl_ln_if_184_acc_nl[14:0];
  assign ln_if_184_acc_itm_14_1 = readslicef_15_1_14(ln_if_184_acc_nl);
  assign nl_ln_if_183_acc_nl = conv_u2u_9_10(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:5])
      + 10'b1111111101;
  assign ln_if_183_acc_nl = nl_ln_if_183_acc_nl[9:0];
  assign ln_if_183_acc_itm_9_1 = readslicef_10_1_9(ln_if_183_acc_nl);
  assign nl_ln_if_182_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110011111;
  assign ln_if_182_acc_nl = nl_ln_if_182_acc_nl[14:0];
  assign ln_if_182_acc_itm_14_1 = readslicef_15_1_14(ln_if_182_acc_nl);
  assign nl_ln_if_181_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111001111;
  assign ln_if_181_acc_nl = nl_ln_if_181_acc_nl[13:0];
  assign ln_if_181_acc_itm_13_1 = readslicef_14_1_13(ln_if_181_acc_nl);
  assign nl_ln_if_180_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110011101;
  assign ln_if_180_acc_nl = nl_ln_if_180_acc_nl[14:0];
  assign ln_if_180_acc_itm_14_1 = readslicef_15_1_14(ln_if_180_acc_nl);
  assign nl_ln_if_179_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111100111;
  assign ln_if_179_acc_nl = nl_ln_if_179_acc_nl[12:0];
  assign ln_if_179_acc_itm_12_1 = readslicef_13_1_12(ln_if_179_acc_nl);
  assign nl_ln_if_178_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110011011;
  assign ln_if_178_acc_nl = nl_ln_if_178_acc_nl[14:0];
  assign ln_if_178_acc_itm_14_1 = readslicef_15_1_14(ln_if_178_acc_nl);
  assign nl_ln_if_177_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111001101;
  assign ln_if_177_acc_nl = nl_ln_if_177_acc_nl[13:0];
  assign ln_if_177_acc_itm_13_1 = readslicef_14_1_13(ln_if_177_acc_nl);
  assign nl_ln_if_176_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110011001;
  assign ln_if_176_acc_nl = nl_ln_if_176_acc_nl[14:0];
  assign ln_if_176_acc_itm_14_1 = readslicef_15_1_14(ln_if_176_acc_nl);
  assign nl_ln_if_175_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:3])
      + 12'b111111110011;
  assign ln_if_175_acc_nl = nl_ln_if_175_acc_nl[11:0];
  assign ln_if_175_acc_itm_11_1 = readslicef_12_1_11(ln_if_175_acc_nl);
  assign nl_ln_if_174_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110010111;
  assign ln_if_174_acc_nl = nl_ln_if_174_acc_nl[14:0];
  assign ln_if_174_acc_itm_14_1 = readslicef_15_1_14(ln_if_174_acc_nl);
  assign nl_ln_if_173_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111001011;
  assign ln_if_173_acc_nl = nl_ln_if_173_acc_nl[13:0];
  assign ln_if_173_acc_itm_13_1 = readslicef_14_1_13(ln_if_173_acc_nl);
  assign nl_ln_if_172_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110010101;
  assign ln_if_172_acc_nl = nl_ln_if_172_acc_nl[14:0];
  assign ln_if_172_acc_itm_14_1 = readslicef_15_1_14(ln_if_172_acc_nl);
  assign nl_ln_if_171_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111100101;
  assign ln_if_171_acc_nl = nl_ln_if_171_acc_nl[12:0];
  assign ln_if_171_acc_itm_12_1 = readslicef_13_1_12(ln_if_171_acc_nl);
  assign nl_ln_if_170_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110010011;
  assign ln_if_170_acc_nl = nl_ln_if_170_acc_nl[14:0];
  assign ln_if_170_acc_itm_14_1 = readslicef_15_1_14(ln_if_170_acc_nl);
  assign nl_ln_if_169_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111001001;
  assign ln_if_169_acc_nl = nl_ln_if_169_acc_nl[13:0];
  assign ln_if_169_acc_itm_13_1 = readslicef_14_1_13(ln_if_169_acc_nl);
  assign nl_ln_if_168_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110010001;
  assign ln_if_168_acc_nl = nl_ln_if_168_acc_nl[14:0];
  assign ln_if_168_acc_itm_14_1 = readslicef_15_1_14(ln_if_168_acc_nl);
  assign nl_ln_if_167_acc_nl = conv_u2u_10_11(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:4])
      + 11'b11111111001;
  assign ln_if_167_acc_nl = nl_ln_if_167_acc_nl[10:0];
  assign ln_if_167_acc_itm_10_1 = readslicef_11_1_10(ln_if_167_acc_nl);
  assign nl_ln_if_166_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110001111;
  assign ln_if_166_acc_nl = nl_ln_if_166_acc_nl[14:0];
  assign ln_if_166_acc_itm_14_1 = readslicef_15_1_14(ln_if_166_acc_nl);
  assign nl_ln_if_165_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111000111;
  assign ln_if_165_acc_nl = nl_ln_if_165_acc_nl[13:0];
  assign ln_if_165_acc_itm_13_1 = readslicef_14_1_13(ln_if_165_acc_nl);
  assign nl_ln_if_164_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110001101;
  assign ln_if_164_acc_nl = nl_ln_if_164_acc_nl[14:0];
  assign ln_if_164_acc_itm_14_1 = readslicef_15_1_14(ln_if_164_acc_nl);
  assign nl_ln_if_163_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111100011;
  assign ln_if_163_acc_nl = nl_ln_if_163_acc_nl[12:0];
  assign ln_if_163_acc_itm_12_1 = readslicef_13_1_12(ln_if_163_acc_nl);
  assign nl_ln_if_162_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110001011;
  assign ln_if_162_acc_nl = nl_ln_if_162_acc_nl[14:0];
  assign ln_if_162_acc_itm_14_1 = readslicef_15_1_14(ln_if_162_acc_nl);
  assign nl_ln_if_161_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111000101;
  assign ln_if_161_acc_nl = nl_ln_if_161_acc_nl[13:0];
  assign ln_if_161_acc_itm_13_1 = readslicef_14_1_13(ln_if_161_acc_nl);
  assign nl_ln_if_160_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110001001;
  assign ln_if_160_acc_nl = nl_ln_if_160_acc_nl[14:0];
  assign ln_if_160_acc_itm_14_1 = readslicef_15_1_14(ln_if_160_acc_nl);
  assign nl_ln_if_159_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:3])
      + 12'b111111110001;
  assign ln_if_159_acc_nl = nl_ln_if_159_acc_nl[11:0];
  assign ln_if_159_acc_itm_11_1 = readslicef_12_1_11(ln_if_159_acc_nl);
  assign nl_ln_if_158_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110000111;
  assign ln_if_158_acc_nl = nl_ln_if_158_acc_nl[14:0];
  assign ln_if_158_acc_itm_14_1 = readslicef_15_1_14(ln_if_158_acc_nl);
  assign nl_ln_if_157_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111000011;
  assign ln_if_157_acc_nl = nl_ln_if_157_acc_nl[13:0];
  assign ln_if_157_acc_itm_13_1 = readslicef_14_1_13(ln_if_157_acc_nl);
  assign nl_ln_if_156_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110000101;
  assign ln_if_156_acc_nl = nl_ln_if_156_acc_nl[14:0];
  assign ln_if_156_acc_itm_14_1 = readslicef_15_1_14(ln_if_156_acc_nl);
  assign nl_ln_if_155_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111100001;
  assign ln_if_155_acc_nl = nl_ln_if_155_acc_nl[12:0];
  assign ln_if_155_acc_itm_12_1 = readslicef_13_1_12(ln_if_155_acc_nl);
  assign nl_ln_if_154_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110000011;
  assign ln_if_154_acc_nl = nl_ln_if_154_acc_nl[14:0];
  assign ln_if_154_acc_itm_14_1 = readslicef_15_1_14(ln_if_154_acc_nl);
  assign nl_ln_if_153_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111111000001;
  assign ln_if_153_acc_nl = nl_ln_if_153_acc_nl[13:0];
  assign ln_if_153_acc_itm_13_1 = readslicef_14_1_13(ln_if_153_acc_nl);
  assign nl_ln_if_152_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111110000001;
  assign ln_if_152_acc_nl = nl_ln_if_152_acc_nl[14:0];
  assign ln_if_152_acc_itm_14_1 = readslicef_15_1_14(ln_if_152_acc_nl);
  assign nl_ln_if_151_acc_nl = conv_u2u_7_8(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:7])
      + 8'b11111111;
  assign ln_if_151_acc_nl = nl_ln_if_151_acc_nl[7:0];
  assign ln_if_151_acc_itm_7_1 = readslicef_8_1_7(ln_if_151_acc_nl);
  assign nl_ln_if_150_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101111111;
  assign ln_if_150_acc_nl = nl_ln_if_150_acc_nl[14:0];
  assign ln_if_150_acc_itm_14_1 = readslicef_15_1_14(ln_if_150_acc_nl);
  assign nl_ln_if_149_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111110111111;
  assign ln_if_149_acc_nl = nl_ln_if_149_acc_nl[13:0];
  assign ln_if_149_acc_itm_13_1 = readslicef_14_1_13(ln_if_149_acc_nl);
  assign nl_ln_if_148_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101111101;
  assign ln_if_148_acc_nl = nl_ln_if_148_acc_nl[14:0];
  assign ln_if_148_acc_itm_14_1 = readslicef_15_1_14(ln_if_148_acc_nl);
  assign nl_ln_if_147_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111011111;
  assign ln_if_147_acc_nl = nl_ln_if_147_acc_nl[12:0];
  assign ln_if_147_acc_itm_12_1 = readslicef_13_1_12(ln_if_147_acc_nl);
  assign nl_ln_if_146_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101111011;
  assign ln_if_146_acc_nl = nl_ln_if_146_acc_nl[14:0];
  assign ln_if_146_acc_itm_14_1 = readslicef_15_1_14(ln_if_146_acc_nl);
  assign nl_ln_if_142_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101110111;
  assign ln_if_142_acc_nl = nl_ln_if_142_acc_nl[14:0];
  assign ln_if_142_acc_itm_14_1 = readslicef_15_1_14(ln_if_142_acc_nl);
  assign nl_ln_if_143_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:3])
      + 12'b111111101111;
  assign ln_if_143_acc_nl = nl_ln_if_143_acc_nl[11:0];
  assign ln_if_143_acc_itm_11_1 = readslicef_12_1_11(ln_if_143_acc_nl);
  assign nl_ln_if_141_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111110111011;
  assign ln_if_141_acc_nl = nl_ln_if_141_acc_nl[13:0];
  assign ln_if_141_acc_itm_13_1 = readslicef_14_1_13(ln_if_141_acc_nl);
  assign nl_ln_if_140_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101110101;
  assign ln_if_140_acc_nl = nl_ln_if_140_acc_nl[14:0];
  assign ln_if_140_acc_itm_14_1 = readslicef_15_1_14(ln_if_140_acc_nl);
  assign nl_ln_if_52_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111010001101;
  assign ln_if_52_acc_nl = nl_ln_if_52_acc_nl[14:0];
  assign ln_if_52_acc_itm_14_1 = readslicef_15_1_14(ln_if_52_acc_nl);
  assign nl_ln_if_53_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111010010001;
  assign ln_if_53_acc_nl = nl_ln_if_53_acc_nl[14:0];
  assign ln_if_53_acc_itm_14_1 = readslicef_15_1_14(ln_if_53_acc_nl);
  assign nl_ln_if_49_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111110100001;
  assign ln_if_49_acc_nl = nl_ln_if_49_acc_nl[12:0];
  assign ln_if_49_acc_itm_12_1 = readslicef_13_1_12(ln_if_49_acc_nl);
  assign nl_ln_if_50_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111010000111;
  assign ln_if_50_acc_nl = nl_ln_if_50_acc_nl[14:0];
  assign ln_if_50_acc_itm_14_1 = readslicef_15_1_14(ln_if_50_acc_nl);
  assign nl_ln_if_6_acc_nl = conv_u2u_8_9(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:6])
      + 9'b111110111;
  assign ln_if_6_acc_nl = nl_ln_if_6_acc_nl[8:0];
  assign ln_if_6_acc_itm_8_1 = readslicef_9_1_8(ln_if_6_acc_nl);
  assign nl_ln_if_7_acc_nl = conv_u2u_5_6(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:9])
      + 6'b111111;
  assign ln_if_7_acc_nl = nl_ln_if_7_acc_nl[5:0];
  assign ln_if_7_acc_itm_5_1 = readslicef_6_1_5(ln_if_7_acc_nl);
  assign nl_ln_if_139_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111011101;
  assign ln_if_139_acc_nl = nl_ln_if_139_acc_nl[12:0];
  assign ln_if_139_acc_itm_12_1 = readslicef_13_1_12(ln_if_139_acc_nl);
  assign nl_ln_if_138_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101110011;
  assign ln_if_138_acc_nl = nl_ln_if_138_acc_nl[14:0];
  assign ln_if_138_acc_itm_14_1 = readslicef_15_1_14(ln_if_138_acc_nl);
  assign nl_ln_if_137_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111110111001;
  assign ln_if_137_acc_nl = nl_ln_if_137_acc_nl[13:0];
  assign ln_if_137_acc_itm_13_1 = readslicef_14_1_13(ln_if_137_acc_nl);
  assign nl_ln_if_136_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101110001;
  assign ln_if_136_acc_nl = nl_ln_if_136_acc_nl[14:0];
  assign ln_if_136_acc_itm_14_1 = readslicef_15_1_14(ln_if_136_acc_nl);
  assign nl_ln_if_135_acc_nl = conv_u2u_10_11(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:4])
      + 11'b11111110111;
  assign ln_if_135_acc_nl = nl_ln_if_135_acc_nl[10:0];
  assign ln_if_135_acc_itm_10_1 = readslicef_11_1_10(ln_if_135_acc_nl);
  assign nl_ln_if_134_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101101111;
  assign ln_if_134_acc_nl = nl_ln_if_134_acc_nl[14:0];
  assign ln_if_134_acc_itm_14_1 = readslicef_15_1_14(ln_if_134_acc_nl);
  assign nl_ln_if_133_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111110110111;
  assign ln_if_133_acc_nl = nl_ln_if_133_acc_nl[13:0];
  assign ln_if_133_acc_itm_13_1 = readslicef_14_1_13(ln_if_133_acc_nl);
  assign nl_ln_if_132_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101101101;
  assign ln_if_132_acc_nl = nl_ln_if_132_acc_nl[14:0];
  assign ln_if_132_acc_itm_14_1 = readslicef_15_1_14(ln_if_132_acc_nl);
  assign nl_ln_if_131_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111011011;
  assign ln_if_131_acc_nl = nl_ln_if_131_acc_nl[12:0];
  assign ln_if_131_acc_itm_12_1 = readslicef_13_1_12(ln_if_131_acc_nl);
  assign nl_ln_if_130_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101101011;
  assign ln_if_130_acc_nl = nl_ln_if_130_acc_nl[14:0];
  assign ln_if_130_acc_itm_14_1 = readslicef_15_1_14(ln_if_130_acc_nl);
  assign nl_ln_if_129_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111110110101;
  assign ln_if_129_acc_nl = nl_ln_if_129_acc_nl[13:0];
  assign ln_if_129_acc_itm_13_1 = readslicef_14_1_13(ln_if_129_acc_nl);
  assign nl_ln_if_128_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101101001;
  assign ln_if_128_acc_nl = nl_ln_if_128_acc_nl[14:0];
  assign ln_if_128_acc_itm_14_1 = readslicef_15_1_14(ln_if_128_acc_nl);
  assign nl_ln_if_127_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:3])
      + 12'b111111101101;
  assign ln_if_127_acc_nl = nl_ln_if_127_acc_nl[11:0];
  assign ln_if_127_acc_itm_11_1 = readslicef_12_1_11(ln_if_127_acc_nl);
  assign nl_ln_if_126_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101100111;
  assign ln_if_126_acc_nl = nl_ln_if_126_acc_nl[14:0];
  assign ln_if_126_acc_itm_14_1 = readslicef_15_1_14(ln_if_126_acc_nl);
  assign nl_ln_if_125_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111110110011;
  assign ln_if_125_acc_nl = nl_ln_if_125_acc_nl[13:0];
  assign ln_if_125_acc_itm_13_1 = readslicef_14_1_13(ln_if_125_acc_nl);
  assign nl_ln_if_124_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101100101;
  assign ln_if_124_acc_nl = nl_ln_if_124_acc_nl[14:0];
  assign ln_if_124_acc_itm_14_1 = readslicef_15_1_14(ln_if_124_acc_nl);
  assign nl_ln_if_123_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111011001;
  assign ln_if_123_acc_nl = nl_ln_if_123_acc_nl[12:0];
  assign ln_if_123_acc_itm_12_1 = readslicef_13_1_12(ln_if_123_acc_nl);
  assign nl_ln_if_122_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101100011;
  assign ln_if_122_acc_nl = nl_ln_if_122_acc_nl[14:0];
  assign ln_if_122_acc_itm_14_1 = readslicef_15_1_14(ln_if_122_acc_nl);
  assign nl_ln_if_121_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111110110001;
  assign ln_if_121_acc_nl = nl_ln_if_121_acc_nl[13:0];
  assign ln_if_121_acc_itm_13_1 = readslicef_14_1_13(ln_if_121_acc_nl);
  assign nl_ln_if_120_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101100001;
  assign ln_if_120_acc_nl = nl_ln_if_120_acc_nl[14:0];
  assign ln_if_120_acc_itm_14_1 = readslicef_15_1_14(ln_if_120_acc_nl);
  assign nl_ln_if_119_acc_nl = conv_u2u_9_10(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:5])
      + 10'b1111111011;
  assign ln_if_119_acc_nl = nl_ln_if_119_acc_nl[9:0];
  assign ln_if_119_acc_itm_9_1 = readslicef_10_1_9(ln_if_119_acc_nl);
  assign nl_ln_if_118_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101011101;
  assign ln_if_118_acc_nl = nl_ln_if_118_acc_nl[14:0];
  assign ln_if_118_acc_itm_14_1 = readslicef_15_1_14(ln_if_118_acc_nl);
  assign nl_ln_if_117_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111110101101;
  assign ln_if_117_acc_nl = nl_ln_if_117_acc_nl[13:0];
  assign ln_if_117_acc_itm_13_1 = readslicef_14_1_13(ln_if_117_acc_nl);
  assign nl_ln_if_116_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101010111;
  assign ln_if_116_acc_nl = nl_ln_if_116_acc_nl[14:0];
  assign ln_if_116_acc_itm_14_1 = readslicef_15_1_14(ln_if_116_acc_nl);
  assign nl_ln_if_115_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101010011;
  assign ln_if_115_acc_nl = nl_ln_if_115_acc_nl[14:0];
  assign ln_if_115_acc_itm_14_1 = readslicef_15_1_14(ln_if_115_acc_nl);
  assign nl_ln_if_114_acc_nl = conv_u2u_10_11(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:4])
      + 11'b11111110101;
  assign ln_if_114_acc_nl = nl_ln_if_114_acc_nl[10:0];
  assign ln_if_114_acc_itm_10_1 = readslicef_11_1_10(ln_if_114_acc_nl);
  assign nl_ln_if_113_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101001101;
  assign ln_if_113_acc_nl = nl_ln_if_113_acc_nl[14:0];
  assign ln_if_113_acc_itm_14_1 = readslicef_15_1_14(ln_if_113_acc_nl);
  assign nl_ln_if_112_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111110100101;
  assign ln_if_112_acc_nl = nl_ln_if_112_acc_nl[13:0];
  assign ln_if_112_acc_itm_13_1 = readslicef_14_1_13(ln_if_112_acc_nl);
  assign nl_ln_if_111_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101000111;
  assign ln_if_111_acc_nl = nl_ln_if_111_acc_nl[14:0];
  assign ln_if_111_acc_itm_14_1 = readslicef_15_1_14(ln_if_111_acc_nl);
  assign nl_ln_if_110_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111010001;
  assign ln_if_110_acc_nl = nl_ln_if_110_acc_nl[12:0];
  assign ln_if_110_acc_itm_12_1 = readslicef_13_1_12(ln_if_110_acc_nl);
  assign nl_ln_if_109_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111101000001;
  assign ln_if_109_acc_nl = nl_ln_if_109_acc_nl[14:0];
  assign ln_if_109_acc_itm_14_1 = readslicef_15_1_14(ln_if_109_acc_nl);
  assign nl_ln_if_108_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111100111101;
  assign ln_if_108_acc_nl = nl_ln_if_108_acc_nl[14:0];
  assign ln_if_108_acc_itm_14_1 = readslicef_15_1_14(ln_if_108_acc_nl);
  assign nl_ln_if_107_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111110011101;
  assign ln_if_107_acc_nl = nl_ln_if_107_acc_nl[13:0];
  assign ln_if_107_acc_itm_13_1 = readslicef_14_1_13(ln_if_107_acc_nl);
  assign nl_ln_if_106_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111100110111;
  assign ln_if_106_acc_nl = nl_ln_if_106_acc_nl[14:0];
  assign ln_if_106_acc_itm_14_1 = readslicef_15_1_14(ln_if_106_acc_nl);
  assign nl_ln_if_105_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111001101;
  assign ln_if_105_acc_nl = nl_ln_if_105_acc_nl[12:0];
  assign ln_if_105_acc_itm_12_1 = readslicef_13_1_12(ln_if_105_acc_nl);
  assign nl_ln_if_104_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111100110001;
  assign ln_if_104_acc_nl = nl_ln_if_104_acc_nl[14:0];
  assign ln_if_104_acc_itm_14_1 = readslicef_15_1_14(ln_if_104_acc_nl);
  assign nl_ln_if_103_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111110010111;
  assign ln_if_103_acc_nl = nl_ln_if_103_acc_nl[13:0];
  assign ln_if_103_acc_itm_13_1 = readslicef_14_1_13(ln_if_103_acc_nl);
  assign nl_ln_if_102_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111100101011;
  assign ln_if_102_acc_nl = nl_ln_if_102_acc_nl[14:0];
  assign ln_if_102_acc_itm_14_1 = readslicef_15_1_14(ln_if_102_acc_nl);
  assign nl_ln_if_101_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111100100111;
  assign ln_if_101_acc_nl = nl_ln_if_101_acc_nl[14:0];
  assign ln_if_101_acc_itm_14_1 = readslicef_15_1_14(ln_if_101_acc_nl);
  assign nl_ln_if_100_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111111001001;
  assign ln_if_100_acc_nl = nl_ln_if_100_acc_nl[12:0];
  assign ln_if_100_acc_itm_12_1 = readslicef_13_1_12(ln_if_100_acc_nl);
  assign nl_ln_if_99_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111100100001;
  assign ln_if_99_acc_nl = nl_ln_if_99_acc_nl[14:0];
  assign ln_if_99_acc_itm_14_1 = readslicef_15_1_14(ln_if_99_acc_nl);
  assign nl_ln_if_98_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111110001111;
  assign ln_if_98_acc_nl = nl_ln_if_98_acc_nl[13:0];
  assign ln_if_98_acc_itm_13_1 = readslicef_14_1_13(ln_if_98_acc_nl);
  assign nl_ln_if_97_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111100011011;
  assign ln_if_97_acc_nl = nl_ln_if_97_acc_nl[14:0];
  assign ln_if_97_acc_itm_14_1 = readslicef_15_1_14(ln_if_97_acc_nl);
  assign nl_ln_if_96_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:3])
      + 12'b111111100011;
  assign ln_if_96_acc_nl = nl_ln_if_96_acc_nl[11:0];
  assign ln_if_96_acc_itm_11_1 = readslicef_12_1_11(ln_if_96_acc_nl);
  assign nl_ln_if_95_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111100010101;
  assign ln_if_95_acc_nl = nl_ln_if_95_acc_nl[14:0];
  assign ln_if_95_acc_itm_14_1 = readslicef_15_1_14(ln_if_95_acc_nl);
  assign nl_ln_if_94_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111100010001;
  assign ln_if_94_acc_nl = nl_ln_if_94_acc_nl[14:0];
  assign ln_if_94_acc_itm_14_1 = readslicef_15_1_14(ln_if_94_acc_nl);
  assign nl_ln_if_93_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111110000111;
  assign ln_if_93_acc_nl = nl_ln_if_93_acc_nl[13:0];
  assign ln_if_93_acc_itm_13_1 = readslicef_14_1_13(ln_if_93_acc_nl);
  assign nl_ln_if_92_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111100001011;
  assign ln_if_92_acc_nl = nl_ln_if_92_acc_nl[14:0];
  assign ln_if_92_acc_itm_14_1 = readslicef_15_1_14(ln_if_92_acc_nl);
  assign nl_ln_if_91_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:3])
      + 12'b111111100001;
  assign ln_if_91_acc_nl = nl_ln_if_91_acc_nl[11:0];
  assign ln_if_91_acc_itm_11_1 = readslicef_12_1_11(ln_if_91_acc_nl);
  assign nl_ln_if_90_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111100000101;
  assign ln_if_90_acc_nl = nl_ln_if_90_acc_nl[14:0];
  assign ln_if_90_acc_itm_14_1 = readslicef_15_1_14(ln_if_90_acc_nl);
  assign nl_ln_if_89_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111110000001;
  assign ln_if_89_acc_nl = nl_ln_if_89_acc_nl[13:0];
  assign ln_if_89_acc_itm_13_1 = readslicef_14_1_13(ln_if_89_acc_nl);
  assign nl_ln_if_88_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111011111111;
  assign ln_if_88_acc_nl = nl_ln_if_88_acc_nl[14:0];
  assign ln_if_88_acc_itm_14_1 = readslicef_15_1_14(ln_if_88_acc_nl);
  assign nl_ln_if_87_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111011111011;
  assign ln_if_87_acc_nl = nl_ln_if_87_acc_nl[14:0];
  assign ln_if_87_acc_itm_14_1 = readslicef_15_1_14(ln_if_87_acc_nl);
  assign nl_ln_if_86_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:3])
      + 12'b111111011111;
  assign ln_if_86_acc_nl = nl_ln_if_86_acc_nl[11:0];
  assign ln_if_86_acc_itm_11_1 = readslicef_12_1_11(ln_if_86_acc_nl);
  assign nl_ln_if_85_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111011110101;
  assign ln_if_85_acc_nl = nl_ln_if_85_acc_nl[14:0];
  assign ln_if_85_acc_itm_14_1 = readslicef_15_1_14(ln_if_85_acc_nl);
  assign nl_ln_if_84_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111101111001;
  assign ln_if_84_acc_nl = nl_ln_if_84_acc_nl[13:0];
  assign ln_if_84_acc_itm_13_1 = readslicef_14_1_13(ln_if_84_acc_nl);
  assign nl_ln_if_83_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111011101111;
  assign ln_if_83_acc_nl = nl_ln_if_83_acc_nl[14:0];
  assign ln_if_83_acc_itm_14_1 = readslicef_15_1_14(ln_if_83_acc_nl);
  assign nl_ln_if_82_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111110111011;
  assign ln_if_82_acc_nl = nl_ln_if_82_acc_nl[12:0];
  assign ln_if_82_acc_itm_12_1 = readslicef_13_1_12(ln_if_82_acc_nl);
  assign nl_ln_if_81_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111011101001;
  assign ln_if_81_acc_nl = nl_ln_if_81_acc_nl[14:0];
  assign ln_if_81_acc_itm_14_1 = readslicef_15_1_14(ln_if_81_acc_nl);
  assign nl_ln_if_80_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111011100101;
  assign ln_if_80_acc_nl = nl_ln_if_80_acc_nl[14:0];
  assign ln_if_80_acc_itm_14_1 = readslicef_15_1_14(ln_if_80_acc_nl);
  assign nl_ln_if_79_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111101110001;
  assign ln_if_79_acc_nl = nl_ln_if_79_acc_nl[13:0];
  assign ln_if_79_acc_itm_13_1 = readslicef_14_1_13(ln_if_79_acc_nl);
  assign nl_ln_if_78_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111011011111;
  assign ln_if_78_acc_nl = nl_ln_if_78_acc_nl[14:0];
  assign ln_if_78_acc_itm_14_1 = readslicef_15_1_14(ln_if_78_acc_nl);
  assign nl_ln_if_77_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111110110111;
  assign ln_if_77_acc_nl = nl_ln_if_77_acc_nl[12:0];
  assign ln_if_77_acc_itm_12_1 = readslicef_13_1_12(ln_if_77_acc_nl);
  assign nl_ln_if_76_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111011011001;
  assign ln_if_76_acc_nl = nl_ln_if_76_acc_nl[14:0];
  assign ln_if_76_acc_itm_14_1 = readslicef_15_1_14(ln_if_76_acc_nl);
  assign nl_ln_if_75_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111101101011;
  assign ln_if_75_acc_nl = nl_ln_if_75_acc_nl[13:0];
  assign ln_if_75_acc_itm_13_1 = readslicef_14_1_13(ln_if_75_acc_nl);
  assign nl_ln_if_74_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111011010011;
  assign ln_if_74_acc_nl = nl_ln_if_74_acc_nl[14:0];
  assign ln_if_74_acc_itm_14_1 = readslicef_15_1_14(ln_if_74_acc_nl);
  assign nl_ln_if_73_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111011001111;
  assign ln_if_73_acc_nl = nl_ln_if_73_acc_nl[14:0];
  assign ln_if_73_acc_itm_14_1 = readslicef_15_1_14(ln_if_73_acc_nl);
  assign nl_ln_if_72_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111110110011;
  assign ln_if_72_acc_nl = nl_ln_if_72_acc_nl[12:0];
  assign ln_if_72_acc_itm_12_1 = readslicef_13_1_12(ln_if_72_acc_nl);
  assign nl_ln_if_71_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111011001001;
  assign ln_if_71_acc_nl = nl_ln_if_71_acc_nl[14:0];
  assign ln_if_71_acc_itm_14_1 = readslicef_15_1_14(ln_if_71_acc_nl);
  assign nl_ln_if_70_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111101100011;
  assign ln_if_70_acc_nl = nl_ln_if_70_acc_nl[13:0];
  assign ln_if_70_acc_itm_13_1 = readslicef_14_1_13(ln_if_70_acc_nl);
  assign nl_ln_if_69_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111011000011;
  assign ln_if_69_acc_nl = nl_ln_if_69_acc_nl[14:0];
  assign ln_if_69_acc_itm_14_1 = readslicef_15_1_14(ln_if_69_acc_nl);
  assign nl_ln_if_68_acc_nl = conv_u2u_8_9(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:6])
      + 9'b111111011;
  assign ln_if_68_acc_nl = nl_ln_if_68_acc_nl[8:0];
  assign ln_if_68_acc_itm_8_1 = readslicef_9_1_8(ln_if_68_acc_nl);
  assign nl_ln_if_67_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111010111101;
  assign ln_if_67_acc_nl = nl_ln_if_67_acc_nl[14:0];
  assign ln_if_67_acc_itm_14_1 = readslicef_15_1_14(ln_if_67_acc_nl);
  assign nl_ln_if_66_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111010111001;
  assign ln_if_66_acc_nl = nl_ln_if_66_acc_nl[14:0];
  assign ln_if_66_acc_itm_14_1 = readslicef_15_1_14(ln_if_66_acc_nl);
  assign nl_ln_if_65_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111101011011;
  assign ln_if_65_acc_nl = nl_ln_if_65_acc_nl[13:0];
  assign ln_if_65_acc_itm_13_1 = readslicef_14_1_13(ln_if_65_acc_nl);
  assign nl_ln_if_64_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111010110011;
  assign ln_if_64_acc_nl = nl_ln_if_64_acc_nl[14:0];
  assign ln_if_64_acc_itm_14_1 = readslicef_15_1_14(ln_if_64_acc_nl);
  assign nl_ln_if_63_acc_nl = conv_u2u_10_11(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:4])
      + 11'b11111101011;
  assign ln_if_63_acc_nl = nl_ln_if_63_acc_nl[10:0];
  assign ln_if_63_acc_itm_10_1 = readslicef_11_1_10(ln_if_63_acc_nl);
  assign nl_ln_if_62_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111010101101;
  assign ln_if_62_acc_nl = nl_ln_if_62_acc_nl[14:0];
  assign ln_if_62_acc_itm_14_1 = readslicef_15_1_14(ln_if_62_acc_nl);
  assign nl_ln_if_61_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111101010101;
  assign ln_if_61_acc_nl = nl_ln_if_61_acc_nl[13:0];
  assign ln_if_61_acc_itm_13_1 = readslicef_14_1_13(ln_if_61_acc_nl);
  assign nl_ln_if_60_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111010100111;
  assign ln_if_60_acc_nl = nl_ln_if_60_acc_nl[14:0];
  assign ln_if_60_acc_itm_14_1 = readslicef_15_1_14(ln_if_60_acc_nl);
  assign nl_ln_if_59_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111010100011;
  assign ln_if_59_acc_nl = nl_ln_if_59_acc_nl[14:0];
  assign ln_if_59_acc_itm_14_1 = readslicef_15_1_14(ln_if_59_acc_nl);
  assign nl_ln_if_58_acc_nl = conv_u2u_9_10(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:5])
      + 10'b1111110101;
  assign ln_if_58_acc_nl = nl_ln_if_58_acc_nl[9:0];
  assign ln_if_58_acc_itm_9_1 = readslicef_10_1_9(ln_if_58_acc_nl);
  assign nl_ln_if_57_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111010011101;
  assign ln_if_57_acc_nl = nl_ln_if_57_acc_nl[14:0];
  assign ln_if_57_acc_itm_14_1 = readslicef_15_1_14(ln_if_57_acc_nl);
  assign nl_ln_if_56_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111101001101;
  assign ln_if_56_acc_nl = nl_ln_if_56_acc_nl[13:0];
  assign ln_if_56_acc_itm_13_1 = readslicef_14_1_13(ln_if_56_acc_nl);
  assign nl_ln_if_55_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111010010111;
  assign ln_if_55_acc_nl = nl_ln_if_55_acc_nl[14:0];
  assign ln_if_55_acc_itm_14_1 = readslicef_15_1_14(ln_if_55_acc_nl);
  assign nl_ln_if_54_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111110100101;
  assign ln_if_54_acc_nl = nl_ln_if_54_acc_nl[12:0];
  assign ln_if_54_acc_itm_12_1 = readslicef_13_1_12(ln_if_54_acc_nl);
  assign nl_ln_if_51_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111101000101;
  assign ln_if_51_acc_nl = nl_ln_if_51_acc_nl[13:0];
  assign ln_if_51_acc_itm_13_1 = readslicef_14_1_13(ln_if_51_acc_nl);
  assign nl_ln_if_48_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111010000001;
  assign ln_if_48_acc_nl = nl_ln_if_48_acc_nl[14:0];
  assign ln_if_48_acc_itm_14_1 = readslicef_15_1_14(ln_if_48_acc_nl);
  assign nl_ln_if_47_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111100111111;
  assign ln_if_47_acc_nl = nl_ln_if_47_acc_nl[13:0];
  assign ln_if_47_acc_itm_13_1 = readslicef_14_1_13(ln_if_47_acc_nl);
  assign nl_ln_if_46_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111001111011;
  assign ln_if_46_acc_nl = nl_ln_if_46_acc_nl[14:0];
  assign ln_if_46_acc_itm_14_1 = readslicef_15_1_14(ln_if_46_acc_nl);
  assign nl_ln_if_45_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111001110111;
  assign ln_if_45_acc_nl = nl_ln_if_45_acc_nl[14:0];
  assign ln_if_45_acc_itm_14_1 = readslicef_15_1_14(ln_if_45_acc_nl);
  assign nl_ln_if_44_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111110011101;
  assign ln_if_44_acc_nl = nl_ln_if_44_acc_nl[12:0];
  assign ln_if_44_acc_itm_12_1 = readslicef_13_1_12(ln_if_44_acc_nl);
  assign nl_ln_if_43_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111001110001;
  assign ln_if_43_acc_nl = nl_ln_if_43_acc_nl[14:0];
  assign ln_if_43_acc_itm_14_1 = readslicef_15_1_14(ln_if_43_acc_nl);
  assign nl_ln_if_42_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111100110111;
  assign ln_if_42_acc_nl = nl_ln_if_42_acc_nl[13:0];
  assign ln_if_42_acc_itm_13_1 = readslicef_14_1_13(ln_if_42_acc_nl);
  assign nl_ln_if_41_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111001101011;
  assign ln_if_41_acc_nl = nl_ln_if_41_acc_nl[14:0];
  assign ln_if_41_acc_itm_14_1 = readslicef_15_1_14(ln_if_41_acc_nl);
  assign nl_ln_if_40_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:3])
      + 12'b111111001101;
  assign ln_if_40_acc_nl = nl_ln_if_40_acc_nl[11:0];
  assign ln_if_40_acc_itm_11_1 = readslicef_12_1_11(ln_if_40_acc_nl);
  assign nl_ln_if_39_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111001100101;
  assign ln_if_39_acc_nl = nl_ln_if_39_acc_nl[14:0];
  assign ln_if_39_acc_itm_14_1 = readslicef_15_1_14(ln_if_39_acc_nl);
  assign nl_ln_if_38_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111001100001;
  assign ln_if_38_acc_nl = nl_ln_if_38_acc_nl[14:0];
  assign ln_if_38_acc_itm_14_1 = readslicef_15_1_14(ln_if_38_acc_nl);
  assign nl_ln_if_37_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111100101111;
  assign ln_if_37_acc_nl = nl_ln_if_37_acc_nl[13:0];
  assign ln_if_37_acc_itm_13_1 = readslicef_14_1_13(ln_if_37_acc_nl);
  assign nl_ln_if_36_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111001011011;
  assign ln_if_36_acc_nl = nl_ln_if_36_acc_nl[14:0];
  assign ln_if_36_acc_itm_14_1 = readslicef_15_1_14(ln_if_36_acc_nl);
  assign nl_ln_if_35_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:3])
      + 12'b111111001011;
  assign ln_if_35_acc_nl = nl_ln_if_35_acc_nl[11:0];
  assign ln_if_35_acc_itm_11_1 = readslicef_12_1_11(ln_if_35_acc_nl);
  assign nl_ln_if_34_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111001010101;
  assign ln_if_34_acc_nl = nl_ln_if_34_acc_nl[14:0];
  assign ln_if_34_acc_itm_14_1 = readslicef_15_1_14(ln_if_34_acc_nl);
  assign nl_ln_if_33_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111100101001;
  assign ln_if_33_acc_nl = nl_ln_if_33_acc_nl[13:0];
  assign ln_if_33_acc_itm_13_1 = readslicef_14_1_13(ln_if_33_acc_nl);
  assign nl_ln_if_32_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111001001111;
  assign ln_if_32_acc_nl = nl_ln_if_32_acc_nl[14:0];
  assign ln_if_32_acc_itm_14_1 = readslicef_15_1_14(ln_if_32_acc_nl);
  assign nl_ln_if_31_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111001001011;
  assign ln_if_31_acc_nl = nl_ln_if_31_acc_nl[14:0];
  assign ln_if_31_acc_itm_14_1 = readslicef_15_1_14(ln_if_31_acc_nl);
  assign nl_ln_if_30_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:3])
      + 12'b111111001001;
  assign ln_if_30_acc_nl = nl_ln_if_30_acc_nl[11:0];
  assign ln_if_30_acc_itm_11_1 = readslicef_12_1_11(ln_if_30_acc_nl);
  assign nl_ln_if_29_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111001000101;
  assign ln_if_29_acc_nl = nl_ln_if_29_acc_nl[14:0];
  assign ln_if_29_acc_itm_14_1 = readslicef_15_1_14(ln_if_29_acc_nl);
  assign nl_ln_if_28_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111100100001;
  assign ln_if_28_acc_nl = nl_ln_if_28_acc_nl[13:0];
  assign ln_if_28_acc_itm_13_1 = readslicef_14_1_13(ln_if_28_acc_nl);
  assign nl_ln_if_27_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111000111111;
  assign ln_if_27_acc_nl = nl_ln_if_27_acc_nl[14:0];
  assign ln_if_27_acc_itm_14_1 = readslicef_15_1_14(ln_if_27_acc_nl);
  assign nl_ln_if_26_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111110001111;
  assign ln_if_26_acc_nl = nl_ln_if_26_acc_nl[12:0];
  assign ln_if_26_acc_itm_12_1 = readslicef_13_1_12(ln_if_26_acc_nl);
  assign nl_ln_if_25_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111000111001;
  assign ln_if_25_acc_nl = nl_ln_if_25_acc_nl[14:0];
  assign ln_if_25_acc_itm_14_1 = readslicef_15_1_14(ln_if_25_acc_nl);
  assign nl_ln_if_24_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111000110101;
  assign ln_if_24_acc_nl = nl_ln_if_24_acc_nl[14:0];
  assign ln_if_24_acc_itm_14_1 = readslicef_15_1_14(ln_if_24_acc_nl);
  assign nl_ln_if_23_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111100011001;
  assign ln_if_23_acc_nl = nl_ln_if_23_acc_nl[13:0];
  assign ln_if_23_acc_itm_13_1 = readslicef_14_1_13(ln_if_23_acc_nl);
  assign nl_ln_if_22_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111000101111;
  assign ln_if_22_acc_nl = nl_ln_if_22_acc_nl[14:0];
  assign ln_if_22_acc_itm_14_1 = readslicef_15_1_14(ln_if_22_acc_nl);
  assign nl_ln_if_21_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111110001011;
  assign ln_if_21_acc_nl = nl_ln_if_21_acc_nl[12:0];
  assign ln_if_21_acc_itm_12_1 = readslicef_13_1_12(ln_if_21_acc_nl);
  assign nl_ln_if_20_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111000101001;
  assign ln_if_20_acc_nl = nl_ln_if_20_acc_nl[14:0];
  assign ln_if_20_acc_itm_14_1 = readslicef_15_1_14(ln_if_20_acc_nl);
  assign nl_ln_if_19_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111100010011;
  assign ln_if_19_acc_nl = nl_ln_if_19_acc_nl[13:0];
  assign ln_if_19_acc_itm_13_1 = readslicef_14_1_13(ln_if_19_acc_nl);
  assign nl_ln_if_18_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111000100011;
  assign ln_if_18_acc_nl = nl_ln_if_18_acc_nl[14:0];
  assign ln_if_18_acc_itm_14_1 = readslicef_15_1_14(ln_if_18_acc_nl);
  assign nl_ln_if_17_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111000011111;
  assign ln_if_17_acc_nl = nl_ln_if_17_acc_nl[14:0];
  assign ln_if_17_acc_itm_14_1 = readslicef_15_1_14(ln_if_17_acc_nl);
  assign nl_ln_if_16_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:2])
      + 13'b1111110000111;
  assign ln_if_16_acc_nl = nl_ln_if_16_acc_nl[12:0];
  assign ln_if_16_acc_itm_12_1 = readslicef_13_1_12(ln_if_16_acc_nl);
  assign nl_ln_if_15_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111000011001;
  assign ln_if_15_acc_nl = nl_ln_if_15_acc_nl[14:0];
  assign ln_if_15_acc_itm_14_1 = readslicef_15_1_14(ln_if_15_acc_nl);
  assign nl_ln_if_14_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111100001011;
  assign ln_if_14_acc_nl = nl_ln_if_14_acc_nl[13:0];
  assign ln_if_14_acc_itm_13_1 = readslicef_14_1_13(ln_if_14_acc_nl);
  assign nl_ln_if_13_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111000010011;
  assign ln_if_13_acc_nl = nl_ln_if_13_acc_nl[14:0];
  assign ln_if_13_acc_itm_14_1 = readslicef_15_1_14(ln_if_13_acc_nl);
  assign nl_ln_if_12_acc_nl = conv_u2u_10_11(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:4])
      + 11'b11111100001;
  assign ln_if_12_acc_nl = nl_ln_if_12_acc_nl[10:0];
  assign ln_if_12_acc_itm_10_1 = readslicef_11_1_10(ln_if_12_acc_nl);
  assign nl_ln_if_11_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111000001101;
  assign ln_if_11_acc_nl = nl_ln_if_11_acc_nl[14:0];
  assign ln_if_11_acc_itm_14_1 = readslicef_15_1_14(ln_if_11_acc_nl);
  assign nl_ln_if_10_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111000001001;
  assign ln_if_10_acc_nl = nl_ln_if_10_acc_nl[14:0];
  assign ln_if_10_acc_itm_14_1 = readslicef_15_1_14(ln_if_10_acc_nl);
  assign nl_ln_if_9_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:1])
      + 14'b11111100000011;
  assign ln_if_9_acc_nl = nl_ln_if_9_acc_nl[13:0];
  assign ln_if_9_acc_itm_13_1 = readslicef_14_1_13(ln_if_9_acc_nl);
  assign nl_ln_if_8_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1)
      + 15'b111111000000011;
  assign ln_if_8_acc_nl = nl_ln_if_8_acc_nl[14:0];
  assign ln_if_8_acc_itm_14_1 = readslicef_15_1_14(ln_if_8_acc_nl);
  assign nl_ln_if_4_acc_nl = conv_u2u_8_9(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:6])
      + 9'b111110101;
  assign ln_if_4_acc_nl = nl_ln_if_4_acc_nl[8:0];
  assign ln_if_4_acc_itm_8_1 = readslicef_9_1_8(ln_if_4_acc_nl);
  assign nl_ln_if_5_acc_nl = conv_u2u_7_8(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:7])
      + 8'b11111011;
  assign ln_if_5_acc_nl = nl_ln_if_5_acc_nl[7:0];
  assign ln_if_5_acc_itm_7_1 = readslicef_8_1_7(ln_if_5_acc_nl);
  assign nl_ln_if_3_acc_nl = conv_u2u_6_7(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:8])
      + 7'b1111101;
  assign ln_if_3_acc_nl = nl_ln_if_3_acc_nl[6:0];
  assign ln_if_3_acc_itm_6_1 = readslicef_7_1_6(ln_if_3_acc_nl);
  assign nl_ln_if_2_acc_nl = conv_u2u_8_9(operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1[13:6])
      + 9'b111110011;
  assign ln_if_2_acc_nl = nl_ln_if_2_acc_nl[8:0];
  assign ln_if_2_acc_itm_8_1 = readslicef_9_1_8(ln_if_2_acc_nl);
  assign if_4_for_and_stg_1_3_sva_1 = (j_1_3_0_lpi_1_dfm_2_0_1[1:0]==2'b11);
  assign if_4_for_and_stg_1_0_sva_1 = ~((j_1_3_0_lpi_1_dfm_2_0_1[1:0]!=2'b00));
  assign if_4_for_and_stg_1_2_sva_1 = (j_1_3_0_lpi_1_dfm_2_0_1[1:0]==2'b10);
  assign if_4_for_and_stg_1_1_sva_1 = (j_1_3_0_lpi_1_dfm_2_0_1[1:0]==2'b01);
  assign ln_1_nor_33_cse_1 = ~((~(ln_1_land_3_lpi_1_dfm_1 | ln_1_land_4_lpi_1_dfm_1
      | ln_1_and_2_ssc_1)) | ln_1_land_6_lpi_1_dfm_1);
  assign ln_1_land_17_lpi_1_dfm_1 = ln_1_if_16_acc_itm_12_1 & (~ ln_1_if_17_acc_itm_14_1);
  assign ln_1_land_18_lpi_1_dfm_1 = ln_1_if_17_acc_itm_14_1 & (~ ln_1_if_18_acc_itm_14_1);
  assign ln_1_land_19_lpi_1_dfm_1 = ln_1_if_18_acc_itm_14_1 & (~ ln_1_if_19_acc_itm_13_1);
  assign ln_1_land_20_lpi_1_dfm_1 = ln_1_if_19_acc_itm_13_1 & (~ ln_1_if_20_acc_itm_14_1);
  assign ln_1_land_21_lpi_1_dfm_1 = ln_1_if_20_acc_itm_14_1 & (~ ln_1_if_21_acc_itm_12_1);
  assign ln_1_land_22_lpi_1_dfm_1 = ln_1_if_21_acc_itm_12_1 & (~ ln_1_if_22_acc_itm_14_1);
  assign ln_1_land_23_lpi_1_dfm_1 = ln_1_if_22_acc_itm_14_1 & (~ ln_1_if_23_acc_itm_13_1);
  assign ln_1_land_24_lpi_1_dfm_1 = ln_1_if_23_acc_itm_13_1 & (~ ln_1_if_24_acc_itm_14_1);
  assign ln_1_land_25_lpi_1_dfm_1 = ln_1_if_24_acc_itm_14_1 & (~ ln_1_if_25_acc_itm_14_1);
  assign ln_1_land_26_lpi_1_dfm_1 = ln_1_if_25_acc_itm_14_1 & (~ ln_1_if_26_acc_itm_12_1);
  assign ln_1_land_27_lpi_1_dfm_1 = ln_1_if_26_acc_itm_12_1 & (~ ln_1_if_27_acc_itm_14_1);
  assign ln_1_land_28_lpi_1_dfm_1 = ln_1_if_27_acc_itm_14_1 & (~ ln_1_if_28_acc_itm_13_1);
  assign ln_1_land_29_lpi_1_dfm_1 = ln_1_if_28_acc_itm_13_1 & (~ ln_1_if_29_acc_itm_14_1);
  assign ln_1_land_30_lpi_1_dfm_1 = ln_1_if_29_acc_itm_14_1 & (~ ln_1_if_30_acc_itm_11_1);
  assign ln_1_land_31_lpi_1_dfm_1 = ln_1_if_30_acc_itm_11_1 & (~ ln_1_if_31_acc_itm_14_1);
  assign ln_1_land_32_lpi_1_dfm_1 = ln_1_if_31_acc_itm_14_1 & (~ ln_1_if_32_acc_itm_14_1);
  assign ln_1_land_33_lpi_1_dfm_1 = ln_1_if_32_acc_itm_14_1 & (~ ln_1_if_33_acc_itm_13_1);
  assign ln_1_land_34_lpi_1_dfm_1 = ln_1_if_33_acc_itm_13_1 & (~ ln_1_if_34_acc_itm_14_1);
  assign ln_1_land_35_lpi_1_dfm_1 = ln_1_if_34_acc_itm_14_1 & (~ ln_1_if_35_acc_itm_11_1);
  assign ln_1_land_36_lpi_1_dfm_1 = ln_1_if_35_acc_itm_11_1 & (~ ln_1_if_36_acc_itm_14_1);
  assign ln_1_land_37_lpi_1_dfm_1 = ln_1_if_36_acc_itm_14_1 & (~ ln_1_if_37_acc_itm_13_1);
  assign ln_1_land_38_lpi_1_dfm_1 = ln_1_if_37_acc_itm_13_1 & (~ ln_1_if_38_acc_itm_14_1);
  assign ln_1_land_39_lpi_1_dfm_1 = ln_1_if_38_acc_itm_14_1 & (~ ln_1_if_39_acc_itm_14_1);
  assign ln_1_land_40_lpi_1_dfm_1 = ln_1_if_39_acc_itm_14_1 & (~ ln_1_if_40_acc_itm_11_1);
  assign ln_1_land_41_lpi_1_dfm_1 = ln_1_if_40_acc_itm_11_1 & (~ ln_1_if_41_acc_itm_14_1);
  assign ln_1_land_42_lpi_1_dfm_1 = ln_1_if_41_acc_itm_14_1 & (~ ln_1_if_42_acc_itm_13_1);
  assign ln_1_land_43_lpi_1_dfm_1 = ln_1_if_42_acc_itm_13_1 & (~ ln_1_if_43_acc_itm_14_1);
  assign ln_1_land_44_lpi_1_dfm_1 = ln_1_if_43_acc_itm_14_1 & (~ ln_1_if_44_acc_itm_12_1);
  assign ln_1_land_45_lpi_1_dfm_1 = ln_1_if_44_acc_itm_12_1 & (~ ln_1_if_45_acc_itm_14_1);
  assign ln_1_land_46_lpi_1_dfm_1 = ln_1_if_45_acc_itm_14_1 & (~ ln_1_if_46_acc_itm_14_1);
  assign ln_1_land_47_lpi_1_dfm_1 = ln_1_if_46_acc_itm_14_1 & (~ ln_1_if_47_acc_itm_13_1);
  assign ln_1_land_48_lpi_1_dfm_1 = ln_1_if_47_acc_itm_13_1 & (~ ln_1_if_48_acc_itm_14_1);
  assign ln_1_land_49_lpi_1_dfm_1 = ln_1_if_48_acc_itm_14_1 & (~ ln_1_if_49_acc_itm_12_1);
  assign ln_1_if_50_ln_1_if_50_and_seb_1 = ln_1_if_49_acc_itm_12_1 & (~ ln_1_if_50_acc_itm_14_1);
  assign ln_1_land_51_lpi_1_dfm_1 = ln_1_if_50_acc_itm_14_1 & (~ ln_1_if_51_acc_itm_13_1);
  assign ln_1_land_52_lpi_1_dfm_1 = ln_1_if_51_acc_itm_13_1 & (~ ln_1_if_52_acc_itm_14_1);
  assign ln_1_land_77_lpi_1_dfm_1 = ln_1_if_76_acc_itm_14_1 & (~ ln_1_if_77_acc_itm_12_1);
  assign ln_1_land_78_lpi_1_dfm_1 = ln_1_if_77_acc_itm_12_1 & (~ ln_1_if_78_acc_itm_14_1);
  assign ln_1_land_79_lpi_1_dfm_1 = ln_1_if_78_acc_itm_14_1 & (~ ln_1_if_79_acc_itm_13_1);
  assign ln_1_land_80_lpi_1_dfm_1 = ln_1_if_79_acc_itm_13_1 & (~ ln_1_if_80_acc_itm_14_1);
  assign ln_1_land_81_lpi_1_dfm_1 = ln_1_if_80_acc_itm_14_1 & (~ ln_1_if_81_acc_itm_14_1);
  assign ln_1_land_82_lpi_1_dfm_1 = ln_1_if_81_acc_itm_14_1 & (~ ln_1_if_82_acc_itm_12_1);
  assign ln_1_land_83_lpi_1_dfm_1 = ln_1_if_82_acc_itm_12_1 & (~ ln_1_if_83_acc_itm_14_1);
  assign ln_1_land_84_lpi_1_dfm_1 = ln_1_if_83_acc_itm_14_1 & (~ ln_1_if_84_acc_itm_13_1);
  assign ln_1_land_85_lpi_1_dfm_1 = ln_1_if_84_acc_itm_13_1 & (~ ln_1_if_85_acc_itm_14_1);
  assign ln_1_land_86_lpi_1_dfm_1 = ln_1_if_85_acc_itm_14_1 & (~ ln_1_if_86_acc_itm_11_1);
  assign ln_1_land_87_lpi_1_dfm_1 = ln_1_if_86_acc_itm_11_1 & (~ ln_1_if_87_acc_itm_14_1);
  assign ln_1_land_88_lpi_1_dfm_1 = ln_1_if_87_acc_itm_14_1 & (~ ln_1_if_88_acc_itm_14_1);
  assign ln_1_land_89_lpi_1_dfm_1 = ln_1_if_88_acc_itm_14_1 & (~ ln_1_if_89_acc_itm_13_1);
  assign ln_1_land_90_lpi_1_dfm_1 = ln_1_if_89_acc_itm_13_1 & (~ ln_1_if_90_acc_itm_14_1);
  assign ln_1_land_91_lpi_1_dfm_1 = ln_1_if_90_acc_itm_14_1 & (~ ln_1_if_91_acc_itm_11_1);
  assign ln_1_land_92_lpi_1_dfm_1 = ln_1_if_91_acc_itm_11_1 & (~ ln_1_if_92_acc_itm_14_1);
  assign ln_1_land_93_lpi_1_dfm_1 = ln_1_if_92_acc_itm_14_1 & (~ ln_1_if_93_acc_itm_13_1);
  assign ln_1_land_94_lpi_1_dfm_1 = ln_1_if_93_acc_itm_13_1 & (~ ln_1_if_94_acc_itm_14_1);
  assign ln_1_land_95_lpi_1_dfm_1 = ln_1_if_94_acc_itm_14_1 & (~ ln_1_if_95_acc_itm_14_1);
  assign ln_1_land_96_lpi_1_dfm_1 = ln_1_if_95_acc_itm_14_1 & (~ ln_1_if_96_acc_itm_11_1);
  assign ln_1_land_97_lpi_1_dfm_1 = ln_1_if_96_acc_itm_11_1 & (~ ln_1_if_97_acc_itm_14_1);
  assign ln_1_land_114_lpi_1_dfm_1 = ln_1_if_113_acc_itm_14_1 & (~ ln_1_if_114_acc_itm_10_1);
  assign ln_1_land_115_lpi_1_dfm_1 = ln_1_if_114_acc_itm_10_1 & (~ ln_1_if_115_acc_itm_14_1);
  assign ln_1_land_116_lpi_1_dfm_1 = ln_1_if_115_acc_itm_14_1 & (~ ln_1_if_116_acc_itm_14_1);
  assign ln_1_land_117_lpi_1_dfm_1 = ln_1_if_116_acc_itm_14_1 & (~ ln_1_if_117_acc_itm_13_1);
  assign ln_1_land_118_lpi_1_dfm_1 = ln_1_if_117_acc_itm_13_1 & (~ ln_1_if_118_acc_itm_14_1);
  assign ln_1_land_119_lpi_1_dfm_1 = ln_1_if_118_acc_itm_14_1 & (~ ln_1_if_119_acc_itm_9_1);
  assign ln_1_land_120_lpi_1_dfm_1 = ln_1_if_119_acc_itm_9_1 & (~ ln_1_if_120_acc_itm_14_1);
  assign ln_1_land_121_lpi_1_dfm_1 = ln_1_if_120_acc_itm_14_1 & (~ ln_1_if_121_acc_itm_13_1);
  assign ln_1_land_122_lpi_1_dfm_1 = ln_1_if_121_acc_itm_13_1 & (~ ln_1_if_122_acc_itm_14_1);
  assign ln_1_land_123_lpi_1_dfm_1 = ln_1_if_122_acc_itm_14_1 & (~ ln_1_if_123_acc_itm_12_1);
  assign ln_1_land_124_lpi_1_dfm_1 = ln_1_if_123_acc_itm_12_1 & (~ ln_1_if_124_acc_itm_14_1);
  assign ln_1_land_125_lpi_1_dfm_1 = ln_1_if_124_acc_itm_14_1 & (~ ln_1_if_125_acc_itm_13_1);
  assign ln_1_land_126_lpi_1_dfm_1 = ln_1_if_125_acc_itm_13_1 & (~ ln_1_if_126_acc_itm_14_1);
  assign ln_1_land_127_lpi_1_dfm_1 = ln_1_if_126_acc_itm_14_1 & (~ ln_1_if_127_acc_itm_11_1);
  assign ln_1_land_128_lpi_1_dfm_1 = ln_1_if_127_acc_itm_11_1 & (~ ln_1_if_128_acc_itm_14_1);
  assign ln_1_land_129_lpi_1_dfm_1 = ln_1_if_128_acc_itm_14_1 & (~ ln_1_if_129_acc_itm_13_1);
  assign ln_1_land_130_lpi_1_dfm_1 = ln_1_if_129_acc_itm_13_1 & (~ ln_1_if_130_acc_itm_14_1);
  assign ln_1_land_131_lpi_1_dfm_1 = ln_1_if_130_acc_itm_14_1 & (~ ln_1_if_131_acc_itm_12_1);
  assign ln_1_land_132_lpi_1_dfm_1 = ln_1_if_131_acc_itm_12_1 & (~ ln_1_if_132_acc_itm_14_1);
  assign ln_1_land_133_lpi_1_dfm_1 = ln_1_if_132_acc_itm_14_1 & (~ ln_1_if_133_acc_itm_13_1);
  assign ln_1_land_134_lpi_1_dfm_1 = ln_1_if_133_acc_itm_13_1 & (~ ln_1_if_134_acc_itm_14_1);
  assign ln_1_land_135_lpi_1_dfm_1 = ln_1_if_134_acc_itm_14_1 & (~ ln_1_if_135_acc_itm_10_1);
  assign ln_1_land_136_lpi_1_dfm_1 = ln_1_if_135_acc_itm_10_1 & (~ ln_1_if_136_acc_itm_14_1);
  assign ln_1_land_137_lpi_1_dfm_1 = ln_1_if_136_acc_itm_14_1 & (~ ln_1_if_137_acc_itm_13_1);
  assign ln_1_land_138_lpi_1_dfm_1 = ln_1_if_137_acc_itm_13_1 & (~ ln_1_if_138_acc_itm_14_1);
  assign ln_1_land_139_lpi_1_dfm_1 = ln_1_if_138_acc_itm_14_1 & (~ ln_1_if_139_acc_itm_12_1);
  assign ln_1_land_140_lpi_1_dfm_1 = ln_1_if_139_acc_itm_12_1 & (~ ln_1_if_140_acc_itm_14_1);
  assign ln_1_and_48_ssc_1 = ln_1_if_52_acc_itm_14_1 & (~ ln_1_if_53_acc_itm_14_1)
      & (~(ln_1_land_55_lpi_1_dfm_1 | ln_1_land_56_lpi_1_dfm_1)) & (~(ln_1_land_57_lpi_1_dfm_1
      | ln_1_land_58_lpi_1_dfm_1)) & (~(ln_1_land_59_lpi_1_dfm_1 | ln_1_land_60_lpi_1_dfm_1))
      & (~(ln_1_land_61_lpi_1_dfm_1 | ln_1_land_62_lpi_1_dfm_1)) & (~(ln_1_land_63_lpi_1_dfm_1
      | ln_1_land_64_lpi_1_dfm_1)) & (~(ln_1_land_65_lpi_1_dfm_1 | ln_1_land_66_lpi_1_dfm_1))
      & (~(ln_1_land_67_lpi_1_dfm_1 | ln_1_land_68_lpi_1_dfm_1)) & (~(ln_1_land_69_lpi_1_dfm_1
      | ln_1_land_70_lpi_1_dfm_1)) & (~(ln_1_land_71_lpi_1_dfm_1 | ln_1_land_72_lpi_1_dfm_1))
      & (~(ln_1_land_73_lpi_1_dfm_1 | ln_1_land_74_lpi_1_dfm_1)) & (~(ln_1_land_75_lpi_1_dfm_1
      | ln_1_land_76_lpi_1_dfm_1)) & (~(ln_1_land_77_lpi_1_dfm_1 | ln_1_land_78_lpi_1_dfm_1))
      & (~(ln_1_land_79_lpi_1_dfm_1 | ln_1_land_80_lpi_1_dfm_1)) & (~(ln_1_land_81_lpi_1_dfm_1
      | ln_1_land_82_lpi_1_dfm_1)) & (~(ln_1_land_83_lpi_1_dfm_1 | ln_1_land_84_lpi_1_dfm_1))
      & (~(ln_1_land_85_lpi_1_dfm_1 | ln_1_land_86_lpi_1_dfm_1)) & (~(ln_1_land_87_lpi_1_dfm_1
      | ln_1_land_88_lpi_1_dfm_1)) & (~(ln_1_land_89_lpi_1_dfm_1 | ln_1_land_90_lpi_1_dfm_1))
      & (~(ln_1_land_91_lpi_1_dfm_1 | ln_1_land_92_lpi_1_dfm_1)) & (~(ln_1_land_93_lpi_1_dfm_1
      | ln_1_land_94_lpi_1_dfm_1)) & (~(ln_1_land_95_lpi_1_dfm_1 | ln_1_land_96_lpi_1_dfm_1))
      & (~(ln_1_land_97_lpi_1_dfm_1 | ln_1_land_98_lpi_1_dfm_1)) & (~(ln_1_land_99_lpi_1_dfm_1
      | ln_1_land_100_lpi_1_dfm_1)) & (~(ln_1_land_101_lpi_1_dfm_1 | ln_1_land_102_lpi_1_dfm_1))
      & (~(ln_1_land_103_lpi_1_dfm_1 | ln_1_land_104_lpi_1_dfm_1)) & (~(ln_1_land_105_lpi_1_dfm_1
      | ln_1_land_106_lpi_1_dfm_1)) & (~(ln_1_land_107_lpi_1_dfm_1 | ln_1_land_108_lpi_1_dfm_1))
      & (~(ln_1_land_109_lpi_1_dfm_1 | ln_1_land_110_lpi_1_dfm_1)) & (~(ln_1_land_111_lpi_1_dfm_1
      | ln_1_land_112_lpi_1_dfm_1)) & (~(ln_1_land_113_lpi_1_dfm_1 | ln_1_land_114_lpi_1_dfm_1))
      & (~(ln_1_land_115_lpi_1_dfm_1 | ln_1_land_116_lpi_1_dfm_1)) & (~(ln_1_land_117_lpi_1_dfm_1
      | ln_1_land_118_lpi_1_dfm_1)) & (~(ln_1_land_119_lpi_1_dfm_1 | ln_1_land_120_lpi_1_dfm_1))
      & (~(ln_1_land_121_lpi_1_dfm_1 | ln_1_land_122_lpi_1_dfm_1)) & (~(ln_1_land_123_lpi_1_dfm_1
      | ln_1_land_124_lpi_1_dfm_1)) & (~(ln_1_land_125_lpi_1_dfm_1 | ln_1_land_126_lpi_1_dfm_1))
      & (~(ln_1_land_127_lpi_1_dfm_1 | ln_1_land_128_lpi_1_dfm_1)) & (~(ln_1_land_129_lpi_1_dfm_1
      | ln_1_land_130_lpi_1_dfm_1)) & (~(ln_1_land_131_lpi_1_dfm_1 | ln_1_land_132_lpi_1_dfm_1))
      & (~(ln_1_land_133_lpi_1_dfm_1 | ln_1_land_134_lpi_1_dfm_1)) & (~(ln_1_land_135_lpi_1_dfm_1
      | ln_1_land_136_lpi_1_dfm_1)) & (~(ln_1_land_137_lpi_1_dfm_1 | ln_1_land_138_lpi_1_dfm_1))
      & (~(ln_1_land_139_lpi_1_dfm_1 | ln_1_land_140_lpi_1_dfm_1));
  assign ln_1_land_54_lpi_1_dfm_1 = ln_1_if_53_acc_itm_14_1 & (~ ln_1_if_54_acc_itm_12_1);
  assign ln_1_land_55_lpi_1_dfm_1 = ln_1_if_54_acc_itm_12_1 & (~ ln_1_if_55_acc_itm_14_1);
  assign ln_1_land_56_lpi_1_dfm_1 = ln_1_if_55_acc_itm_14_1 & (~ ln_1_if_56_acc_itm_13_1);
  assign ln_1_land_57_lpi_1_dfm_1 = ln_1_if_56_acc_itm_13_1 & (~ ln_1_if_57_acc_itm_14_1);
  assign ln_1_land_58_lpi_1_dfm_1 = ln_1_if_57_acc_itm_14_1 & (~ ln_1_if_58_acc_itm_9_1);
  assign ln_1_land_59_lpi_1_dfm_1 = ln_1_if_58_acc_itm_9_1 & (~ ln_1_if_59_acc_itm_14_1);
  assign ln_1_land_60_lpi_1_dfm_1 = ln_1_if_59_acc_itm_14_1 & (~ ln_1_if_60_acc_itm_14_1);
  assign ln_1_land_61_lpi_1_dfm_1 = ln_1_if_60_acc_itm_14_1 & (~ ln_1_if_61_acc_itm_13_1);
  assign ln_1_land_62_lpi_1_dfm_1 = ln_1_if_61_acc_itm_13_1 & (~ ln_1_if_62_acc_itm_14_1);
  assign ln_1_land_63_lpi_1_dfm_1 = ln_1_if_62_acc_itm_14_1 & (~ ln_1_if_63_acc_itm_10_1);
  assign ln_1_land_64_lpi_1_dfm_1 = ln_1_if_63_acc_itm_10_1 & (~ ln_1_if_64_acc_itm_14_1);
  assign ln_1_land_65_lpi_1_dfm_1 = ln_1_if_64_acc_itm_14_1 & (~ ln_1_if_65_acc_itm_13_1);
  assign ln_1_land_66_lpi_1_dfm_1 = ln_1_if_65_acc_itm_13_1 & (~ ln_1_if_66_acc_itm_14_1);
  assign ln_1_land_67_lpi_1_dfm_1 = ln_1_if_66_acc_itm_14_1 & (~ ln_1_if_67_acc_itm_14_1);
  assign ln_1_land_68_lpi_1_dfm_1 = ln_1_if_67_acc_itm_14_1 & (~ ln_1_if_68_acc_itm_8_1);
  assign ln_1_land_69_lpi_1_dfm_1 = ln_1_if_68_acc_itm_8_1 & (~ ln_1_if_69_acc_itm_14_1);
  assign ln_1_land_70_lpi_1_dfm_1 = ln_1_if_69_acc_itm_14_1 & (~ ln_1_if_70_acc_itm_13_1);
  assign ln_1_land_71_lpi_1_dfm_1 = ln_1_if_70_acc_itm_13_1 & (~ ln_1_if_71_acc_itm_14_1);
  assign ln_1_land_72_lpi_1_dfm_1 = ln_1_if_71_acc_itm_14_1 & (~ ln_1_if_72_acc_itm_12_1);
  assign ln_1_land_73_lpi_1_dfm_1 = ln_1_if_72_acc_itm_12_1 & (~ ln_1_if_73_acc_itm_14_1);
  assign ln_1_land_74_lpi_1_dfm_1 = ln_1_if_73_acc_itm_14_1 & (~ ln_1_if_74_acc_itm_14_1);
  assign ln_1_land_75_lpi_1_dfm_1 = ln_1_if_74_acc_itm_14_1 & (~ ln_1_if_75_acc_itm_13_1);
  assign ln_1_land_76_lpi_1_dfm_1 = ln_1_if_75_acc_itm_13_1 & (~ ln_1_if_76_acc_itm_14_1);
  assign ln_1_land_98_lpi_1_dfm_1 = ln_1_if_97_acc_itm_14_1 & (~ ln_1_if_98_acc_itm_13_1);
  assign ln_1_land_99_lpi_1_dfm_1 = ln_1_if_98_acc_itm_13_1 & (~ ln_1_if_99_acc_itm_14_1);
  assign ln_1_land_100_lpi_1_dfm_1 = ln_1_if_99_acc_itm_14_1 & (~ ln_1_if_100_acc_itm_12_1);
  assign ln_1_land_101_lpi_1_dfm_1 = ln_1_if_100_acc_itm_12_1 & (~ ln_1_if_101_acc_itm_14_1);
  assign ln_1_land_102_lpi_1_dfm_1 = ln_1_if_101_acc_itm_14_1 & (~ ln_1_if_102_acc_itm_14_1);
  assign ln_1_land_103_lpi_1_dfm_1 = ln_1_if_102_acc_itm_14_1 & (~ ln_1_if_103_acc_itm_13_1);
  assign ln_1_land_104_lpi_1_dfm_1 = ln_1_if_103_acc_itm_13_1 & (~ ln_1_if_104_acc_itm_14_1);
  assign ln_1_land_105_lpi_1_dfm_1 = ln_1_if_104_acc_itm_14_1 & (~ ln_1_if_105_acc_itm_12_1);
  assign ln_1_land_106_lpi_1_dfm_1 = ln_1_if_105_acc_itm_12_1 & (~ ln_1_if_106_acc_itm_14_1);
  assign ln_1_land_107_lpi_1_dfm_1 = ln_1_if_106_acc_itm_14_1 & (~ ln_1_if_107_acc_itm_13_1);
  assign ln_1_land_108_lpi_1_dfm_1 = ln_1_if_107_acc_itm_13_1 & (~ ln_1_if_108_acc_itm_14_1);
  assign ln_1_land_109_lpi_1_dfm_1 = ln_1_if_108_acc_itm_14_1 & (~ ln_1_if_109_acc_itm_14_1);
  assign ln_1_land_110_lpi_1_dfm_1 = ln_1_if_109_acc_itm_14_1 & (~ ln_1_if_110_acc_itm_12_1);
  assign ln_1_land_111_lpi_1_dfm_1 = ln_1_if_110_acc_itm_12_1 & (~ ln_1_if_111_acc_itm_14_1);
  assign ln_1_land_112_lpi_1_dfm_1 = ln_1_if_111_acc_itm_14_1 & (~ ln_1_if_112_acc_itm_13_1);
  assign ln_1_land_113_lpi_1_dfm_1 = ln_1_if_112_acc_itm_13_1 & (~ ln_1_if_113_acc_itm_14_1);
  assign ln_1_land_141_lpi_1_dfm_1 = ln_1_if_140_acc_itm_14_1 & (~ ln_1_if_141_acc_itm_13_1);
  assign ln_1_land_142_lpi_1_dfm_1 = ln_1_if_141_acc_itm_13_1 & (~ ln_1_if_142_acc_itm_14_1);
  assign ln_1_and_138_ssc_1 = ln_1_if_142_acc_itm_14_1 & (~ ln_1_if_143_acc_itm_11_1);
  assign ln_1_land_144_lpi_1_dfm_1 = ln_1_if_143_acc_itm_11_1 & (~ ln_1_if_144_acc_itm_14_1);
  assign ln_1_land_172_lpi_1_dfm_1 = ln_1_if_171_acc_itm_12_1 & (~ ln_1_if_172_acc_itm_14_1);
  assign ln_1_land_173_lpi_1_dfm_1 = ln_1_if_172_acc_itm_14_1 & (~ ln_1_if_173_acc_itm_13_1);
  assign ln_1_land_174_lpi_1_dfm_1 = ln_1_if_173_acc_itm_13_1 & (~ ln_1_if_174_acc_itm_14_1);
  assign ln_1_land_175_lpi_1_dfm_1 = ln_1_if_174_acc_itm_14_1 & (~ ln_1_if_175_acc_itm_11_1);
  assign ln_1_land_176_lpi_1_dfm_1 = ln_1_if_175_acc_itm_11_1 & (~ ln_1_if_176_acc_itm_14_1);
  assign ln_1_land_177_lpi_1_dfm_1 = ln_1_if_176_acc_itm_14_1 & (~ ln_1_if_177_acc_itm_13_1);
  assign ln_1_land_178_lpi_1_dfm_1 = ln_1_if_177_acc_itm_13_1 & (~ ln_1_if_178_acc_itm_14_1);
  assign ln_1_land_179_lpi_1_dfm_1 = ln_1_if_178_acc_itm_14_1 & (~ ln_1_if_179_acc_itm_12_1);
  assign ln_1_land_180_lpi_1_dfm_1 = ln_1_if_179_acc_itm_12_1 & (~ ln_1_if_180_acc_itm_14_1);
  assign ln_1_land_181_lpi_1_dfm_1 = ln_1_if_180_acc_itm_14_1 & (~ ln_1_if_181_acc_itm_13_1);
  assign ln_1_land_182_lpi_1_dfm_1 = ln_1_if_181_acc_itm_13_1 & (~ ln_1_if_182_acc_itm_14_1);
  assign ln_1_land_183_lpi_1_dfm_1 = ln_1_if_182_acc_itm_14_1 & (~ ln_1_if_183_acc_itm_9_1);
  assign ln_1_land_184_lpi_1_dfm_1 = ln_1_if_183_acc_itm_9_1 & (~ ln_1_if_184_acc_itm_14_1);
  assign ln_1_land_185_lpi_1_dfm_1 = ln_1_if_184_acc_itm_14_1 & (~ ln_1_if_185_acc_itm_13_1);
  assign ln_1_land_186_lpi_1_dfm_1 = ln_1_if_185_acc_itm_13_1 & (~ ln_1_if_186_acc_itm_14_1);
  assign ln_1_land_187_lpi_1_dfm_1 = ln_1_if_186_acc_itm_14_1 & (~ ln_1_if_187_acc_itm_12_1);
  assign ln_1_land_188_lpi_1_dfm_1 = ln_1_if_187_acc_itm_12_1 & (~ ln_1_if_188_acc_itm_14_1);
  assign ln_1_land_189_lpi_1_dfm_1 = ln_1_if_188_acc_itm_14_1 & (~ ln_1_if_189_acc_itm_13_1);
  assign ln_1_land_190_lpi_1_dfm_1 = ln_1_if_189_acc_itm_13_1 & (~ ln_1_if_190_acc_itm_14_1);
  assign ln_1_land_191_lpi_1_dfm_1 = ln_1_if_190_acc_itm_14_1 & (~ ln_1_if_191_acc_itm_11_1);
  assign ln_1_land_192_lpi_1_dfm_1 = ln_1_if_191_acc_itm_11_1 & (~ ln_1_if_192_acc_itm_14_1);
  assign ln_1_land_193_lpi_1_dfm_1 = ln_1_if_192_acc_itm_14_1 & (~ ln_1_if_193_acc_itm_13_1);
  assign ln_1_land_194_lpi_1_dfm_1 = ln_1_if_193_acc_itm_13_1 & (~ ln_1_if_194_acc_itm_14_1);
  assign ln_1_land_214_lpi_1_dfm_1 = ln_1_if_213_acc_itm_13_1 & (~ ln_1_if_214_acc_itm_14_1);
  assign ln_1_land_215_lpi_1_dfm_1 = ln_1_if_214_acc_itm_14_1 & (~ ln_1_if_215_acc_itm_8_1);
  assign ln_1_land_216_lpi_1_dfm_1 = ln_1_if_215_acc_itm_8_1 & (~ ln_1_if_216_acc_itm_14_1);
  assign ln_1_land_217_lpi_1_dfm_1 = ln_1_if_216_acc_itm_14_1 & (~ ln_1_if_217_acc_itm_13_1);
  assign ln_1_land_218_lpi_1_dfm_1 = ln_1_if_217_acc_itm_13_1 & (~ ln_1_if_218_acc_itm_14_1);
  assign ln_1_land_219_lpi_1_dfm_1 = ln_1_if_218_acc_itm_14_1 & (~ ln_1_if_219_acc_itm_12_1);
  assign ln_1_land_220_lpi_1_dfm_1 = ln_1_if_219_acc_itm_12_1 & (~ ln_1_if_220_acc_itm_14_1);
  assign ln_1_land_221_lpi_1_dfm_1 = ln_1_if_220_acc_itm_14_1 & (~ ln_1_if_221_acc_itm_13_1);
  assign ln_1_land_222_lpi_1_dfm_1 = ln_1_if_221_acc_itm_13_1 & (~ ln_1_if_222_acc_itm_14_1);
  assign ln_1_land_223_lpi_1_dfm_1 = ln_1_if_222_acc_itm_14_1 & (~ ln_1_if_223_acc_itm_11_1);
  assign ln_1_land_224_lpi_1_dfm_1 = ln_1_if_223_acc_itm_11_1 & (~ ln_1_if_224_acc_itm_14_1);
  assign ln_1_land_225_lpi_1_dfm_1 = ln_1_if_224_acc_itm_14_1 & (~ ln_1_if_225_acc_itm_13_1);
  assign ln_1_land_226_lpi_1_dfm_1 = ln_1_if_225_acc_itm_13_1 & (~ ln_1_if_226_acc_itm_14_1);
  assign ln_1_land_227_lpi_1_dfm_1 = ln_1_if_226_acc_itm_14_1 & (~ ln_1_if_227_acc_itm_12_1);
  assign ln_1_land_228_lpi_1_dfm_1 = ln_1_if_227_acc_itm_12_1 & (~ ln_1_if_228_acc_itm_14_1);
  assign ln_1_land_240_lpi_1_dfm_1 = ln_1_if_239_acc_itm_11_1 & (~ ln_1_if_240_acc_itm_14_1);
  assign ln_1_land_241_lpi_1_dfm_1 = ln_1_if_240_acc_itm_14_1 & (~ ln_1_if_241_acc_itm_13_1);
  assign ln_1_land_242_lpi_1_dfm_1 = ln_1_if_241_acc_itm_13_1 & (~ ln_1_if_242_acc_itm_14_1);
  assign ln_1_land_243_lpi_1_dfm_1 = ln_1_if_242_acc_itm_14_1 & (~ ln_1_if_243_acc_itm_12_1);
  assign ln_1_land_244_lpi_1_dfm_1 = ln_1_if_243_acc_itm_12_1 & (~ ln_1_if_244_acc_itm_14_1);
  assign ln_1_and_140_ssc_1 = ln_1_if_144_acc_itm_14_1 & (~ ln_1_if_145_acc_itm_13_1)
      & (~(ln_1_land_147_lpi_1_dfm_1 | ln_1_land_148_lpi_1_dfm_1)) & (~(ln_1_land_149_lpi_1_dfm_1
      | ln_1_land_150_lpi_1_dfm_1)) & (~(ln_1_land_151_lpi_1_dfm_1 | ln_1_land_152_lpi_1_dfm_1))
      & (~(ln_1_land_153_lpi_1_dfm_1 | ln_1_land_154_lpi_1_dfm_1)) & (~(ln_1_land_155_lpi_1_dfm_1
      | ln_1_land_156_lpi_1_dfm_1)) & (~(ln_1_land_157_lpi_1_dfm_1 | ln_1_land_158_lpi_1_dfm_1))
      & (~(ln_1_land_159_lpi_1_dfm_1 | ln_1_land_160_lpi_1_dfm_1)) & (~(ln_1_land_161_lpi_1_dfm_1
      | ln_1_land_162_lpi_1_dfm_1)) & (~(ln_1_land_163_lpi_1_dfm_1 | ln_1_land_164_lpi_1_dfm_1))
      & (~(ln_1_land_165_lpi_1_dfm_1 | ln_1_land_166_lpi_1_dfm_1)) & (~(ln_1_land_167_lpi_1_dfm_1
      | ln_1_land_168_lpi_1_dfm_1)) & (~(ln_1_land_169_lpi_1_dfm_1 | ln_1_land_170_lpi_1_dfm_1))
      & (~(ln_1_land_171_lpi_1_dfm_1 | ln_1_land_172_lpi_1_dfm_1)) & (~(ln_1_land_173_lpi_1_dfm_1
      | ln_1_land_174_lpi_1_dfm_1)) & (~(ln_1_land_175_lpi_1_dfm_1 | ln_1_land_176_lpi_1_dfm_1))
      & (~(ln_1_land_177_lpi_1_dfm_1 | ln_1_land_178_lpi_1_dfm_1)) & (~(ln_1_land_179_lpi_1_dfm_1
      | ln_1_land_180_lpi_1_dfm_1)) & (~(ln_1_land_181_lpi_1_dfm_1 | ln_1_land_182_lpi_1_dfm_1))
      & (~(ln_1_land_183_lpi_1_dfm_1 | ln_1_land_184_lpi_1_dfm_1)) & (~(ln_1_land_185_lpi_1_dfm_1
      | ln_1_land_186_lpi_1_dfm_1)) & (~(ln_1_land_187_lpi_1_dfm_1 | ln_1_land_188_lpi_1_dfm_1))
      & (~(ln_1_land_189_lpi_1_dfm_1 | ln_1_land_190_lpi_1_dfm_1)) & (~(ln_1_land_191_lpi_1_dfm_1
      | ln_1_land_192_lpi_1_dfm_1)) & (~(ln_1_land_193_lpi_1_dfm_1 | ln_1_land_194_lpi_1_dfm_1))
      & (~(ln_1_land_195_lpi_1_dfm_1 | ln_1_land_196_lpi_1_dfm_1)) & (~(ln_1_land_197_lpi_1_dfm_1
      | ln_1_land_198_lpi_1_dfm_1)) & (~(ln_1_land_199_lpi_1_dfm_1 | ln_1_land_200_lpi_1_dfm_1))
      & (~(ln_1_land_201_lpi_1_dfm_1 | ln_1_land_202_lpi_1_dfm_1)) & (~(ln_1_land_203_lpi_1_dfm_1
      | ln_1_land_204_lpi_1_dfm_1)) & (~(ln_1_land_205_lpi_1_dfm_1 | ln_1_land_206_lpi_1_dfm_1))
      & (~(ln_1_land_207_lpi_1_dfm_1 | ln_1_land_208_lpi_1_dfm_1)) & (~(ln_1_land_209_lpi_1_dfm_1
      | ln_1_land_210_lpi_1_dfm_1)) & (~(ln_1_land_211_lpi_1_dfm_1 | ln_1_land_212_lpi_1_dfm_1))
      & (~(ln_1_land_213_lpi_1_dfm_1 | ln_1_land_214_lpi_1_dfm_1)) & (~(ln_1_land_215_lpi_1_dfm_1
      | ln_1_land_216_lpi_1_dfm_1)) & (~(ln_1_land_217_lpi_1_dfm_1 | ln_1_land_218_lpi_1_dfm_1))
      & (~(ln_1_land_219_lpi_1_dfm_1 | ln_1_land_220_lpi_1_dfm_1)) & (~(ln_1_land_221_lpi_1_dfm_1
      | ln_1_land_222_lpi_1_dfm_1)) & (~(ln_1_land_223_lpi_1_dfm_1 | ln_1_land_224_lpi_1_dfm_1))
      & (~(ln_1_land_225_lpi_1_dfm_1 | ln_1_land_226_lpi_1_dfm_1)) & (~(ln_1_land_227_lpi_1_dfm_1
      | ln_1_land_228_lpi_1_dfm_1)) & ln_1_and_368_m1c_1;
  assign ln_1_land_146_lpi_1_dfm_1 = ln_1_if_145_acc_itm_13_1 & (~ ln_1_if_146_acc_itm_14_1);
  assign ln_1_land_147_lpi_1_dfm_1 = ln_1_if_146_acc_itm_14_1 & (~ ln_1_if_147_acc_itm_12_1);
  assign ln_1_land_148_lpi_1_dfm_1 = ln_1_if_147_acc_itm_12_1 & (~ ln_1_if_148_acc_itm_14_1);
  assign ln_1_land_149_lpi_1_dfm_1 = ln_1_if_148_acc_itm_14_1 & (~ ln_1_if_149_acc_itm_13_1);
  assign ln_1_land_150_lpi_1_dfm_1 = ln_1_if_149_acc_itm_13_1 & (~ ln_1_if_150_acc_itm_14_1);
  assign ln_1_land_151_lpi_1_dfm_1 = ln_1_if_150_acc_itm_14_1 & (~ ln_1_if_151_acc_itm_7_1);
  assign ln_1_land_152_lpi_1_dfm_1 = ln_1_if_151_acc_itm_7_1 & (~ ln_1_if_152_acc_itm_14_1);
  assign ln_1_land_153_lpi_1_dfm_1 = ln_1_if_152_acc_itm_14_1 & (~ ln_1_if_153_acc_itm_13_1);
  assign ln_1_land_154_lpi_1_dfm_1 = ln_1_if_153_acc_itm_13_1 & (~ ln_1_if_154_acc_itm_14_1);
  assign ln_1_land_155_lpi_1_dfm_1 = ln_1_if_154_acc_itm_14_1 & (~ ln_1_if_155_acc_itm_12_1);
  assign ln_1_land_156_lpi_1_dfm_1 = ln_1_if_155_acc_itm_12_1 & (~ ln_1_if_156_acc_itm_14_1);
  assign ln_1_land_157_lpi_1_dfm_1 = ln_1_if_156_acc_itm_14_1 & (~ ln_1_if_157_acc_itm_13_1);
  assign ln_1_land_158_lpi_1_dfm_1 = ln_1_if_157_acc_itm_13_1 & (~ ln_1_if_158_acc_itm_14_1);
  assign ln_1_land_159_lpi_1_dfm_1 = ln_1_if_158_acc_itm_14_1 & (~ ln_1_if_159_acc_itm_11_1);
  assign ln_1_land_160_lpi_1_dfm_1 = ln_1_if_159_acc_itm_11_1 & (~ ln_1_if_160_acc_itm_14_1);
  assign ln_1_land_161_lpi_1_dfm_1 = ln_1_if_160_acc_itm_14_1 & (~ ln_1_if_161_acc_itm_13_1);
  assign ln_1_land_162_lpi_1_dfm_1 = ln_1_if_161_acc_itm_13_1 & (~ ln_1_if_162_acc_itm_14_1);
  assign ln_1_land_163_lpi_1_dfm_1 = ln_1_if_162_acc_itm_14_1 & (~ ln_1_if_163_acc_itm_12_1);
  assign ln_1_land_164_lpi_1_dfm_1 = ln_1_if_163_acc_itm_12_1 & (~ ln_1_if_164_acc_itm_14_1);
  assign ln_1_land_165_lpi_1_dfm_1 = ln_1_if_164_acc_itm_14_1 & (~ ln_1_if_165_acc_itm_13_1);
  assign ln_1_land_166_lpi_1_dfm_1 = ln_1_if_165_acc_itm_13_1 & (~ ln_1_if_166_acc_itm_14_1);
  assign ln_1_land_167_lpi_1_dfm_1 = ln_1_if_166_acc_itm_14_1 & (~ ln_1_if_167_acc_itm_10_1);
  assign ln_1_land_168_lpi_1_dfm_1 = ln_1_if_167_acc_itm_10_1 & (~ ln_1_if_168_acc_itm_14_1);
  assign ln_1_land_169_lpi_1_dfm_1 = ln_1_if_168_acc_itm_14_1 & (~ ln_1_if_169_acc_itm_13_1);
  assign ln_1_land_170_lpi_1_dfm_1 = ln_1_if_169_acc_itm_13_1 & (~ ln_1_if_170_acc_itm_14_1);
  assign ln_1_land_171_lpi_1_dfm_1 = ln_1_if_170_acc_itm_14_1 & (~ ln_1_if_171_acc_itm_12_1);
  assign ln_1_land_195_lpi_1_dfm_1 = ln_1_if_194_acc_itm_14_1 & (~ ln_1_if_195_acc_itm_12_1);
  assign ln_1_land_196_lpi_1_dfm_1 = ln_1_if_195_acc_itm_12_1 & (~ ln_1_if_196_acc_itm_14_1);
  assign ln_1_land_197_lpi_1_dfm_1 = ln_1_if_196_acc_itm_14_1 & (~ ln_1_if_197_acc_itm_13_1);
  assign ln_1_land_198_lpi_1_dfm_1 = ln_1_if_197_acc_itm_13_1 & (~ ln_1_if_198_acc_itm_14_1);
  assign ln_1_land_199_lpi_1_dfm_1 = ln_1_if_198_acc_itm_14_1 & (~ ln_1_if_199_acc_itm_10_1);
  assign ln_1_land_200_lpi_1_dfm_1 = ln_1_if_199_acc_itm_10_1 & (~ ln_1_if_200_acc_itm_14_1);
  assign ln_1_land_201_lpi_1_dfm_1 = ln_1_if_200_acc_itm_14_1 & (~ ln_1_if_201_acc_itm_13_1);
  assign ln_1_land_202_lpi_1_dfm_1 = ln_1_if_201_acc_itm_13_1 & (~ ln_1_if_202_acc_itm_14_1);
  assign ln_1_land_203_lpi_1_dfm_1 = ln_1_if_202_acc_itm_14_1 & (~ ln_1_if_203_acc_itm_12_1);
  assign ln_1_land_204_lpi_1_dfm_1 = ln_1_if_203_acc_itm_12_1 & (~ ln_1_if_204_acc_itm_14_1);
  assign ln_1_land_205_lpi_1_dfm_1 = ln_1_if_204_acc_itm_14_1 & (~ ln_1_if_205_acc_itm_13_1);
  assign ln_1_land_206_lpi_1_dfm_1 = ln_1_if_205_acc_itm_13_1 & (~ ln_1_if_206_acc_itm_14_1);
  assign ln_1_land_207_lpi_1_dfm_1 = ln_1_if_206_acc_itm_14_1 & (~ ln_1_if_207_acc_itm_11_1);
  assign ln_1_land_208_lpi_1_dfm_1 = ln_1_if_207_acc_itm_11_1 & (~ ln_1_if_208_acc_itm_14_1);
  assign ln_1_land_209_lpi_1_dfm_1 = ln_1_if_208_acc_itm_14_1 & (~ ln_1_if_209_acc_itm_13_1);
  assign ln_1_land_210_lpi_1_dfm_1 = ln_1_if_209_acc_itm_13_1 & (~ ln_1_if_210_acc_itm_14_1);
  assign ln_1_land_211_lpi_1_dfm_1 = ln_1_if_210_acc_itm_14_1 & (~ ln_1_if_211_acc_itm_12_1);
  assign ln_1_land_212_lpi_1_dfm_1 = ln_1_if_211_acc_itm_12_1 & (~ ln_1_if_212_acc_itm_14_1);
  assign ln_1_land_213_lpi_1_dfm_1 = ln_1_if_212_acc_itm_14_1 & (~ ln_1_if_213_acc_itm_13_1);
  assign ln_1_land_229_lpi_1_dfm_1 = ln_1_if_228_acc_itm_14_1 & (~ ln_1_if_229_acc_itm_13_1);
  assign ln_1_land_230_lpi_1_dfm_1 = ln_1_if_229_acc_itm_13_1 & (~ ln_1_if_230_acc_itm_14_1);
  assign ln_1_land_231_lpi_1_dfm_1 = ln_1_if_230_acc_itm_14_1 & (~ ln_1_if_231_acc_itm_10_1);
  assign ln_1_land_232_lpi_1_dfm_1 = ln_1_if_231_acc_itm_10_1 & (~ ln_1_if_232_acc_itm_14_1);
  assign ln_1_land_233_lpi_1_dfm_1 = ln_1_if_232_acc_itm_14_1 & (~ ln_1_if_233_acc_itm_13_1);
  assign ln_1_land_234_lpi_1_dfm_1 = ln_1_if_233_acc_itm_13_1 & (~ ln_1_if_234_acc_itm_14_1);
  assign ln_1_land_235_lpi_1_dfm_1 = ln_1_if_234_acc_itm_14_1 & (~ ln_1_if_235_acc_itm_12_1);
  assign ln_1_land_236_lpi_1_dfm_1 = ln_1_if_235_acc_itm_12_1 & (~ ln_1_if_236_acc_itm_14_1);
  assign ln_1_land_237_lpi_1_dfm_1 = ln_1_if_236_acc_itm_14_1 & (~ ln_1_if_237_acc_itm_13_1);
  assign ln_1_land_238_lpi_1_dfm_1 = ln_1_if_237_acc_itm_13_1 & (~ ln_1_if_238_acc_itm_14_1);
  assign ln_1_land_239_lpi_1_dfm_1 = ln_1_if_238_acc_itm_14_1 & (~ ln_1_if_239_acc_itm_11_1);
  assign nl_ln_1_if_252_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111111101;
  assign ln_1_if_252_acc_nl = nl_ln_1_if_252_acc_nl[12:0];
  assign ln_1_if_252_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_252_acc_nl);
  assign nl_ln_1_if_244_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111111011101;
  assign ln_1_if_244_acc_nl = nl_ln_1_if_244_acc_nl[14:0];
  assign ln_1_if_244_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_244_acc_nl);
  assign nl_ln_1_if_245_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111101111;
  assign ln_1_if_245_acc_nl = nl_ln_1_if_245_acc_nl[13:0];
  assign ln_1_if_245_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_245_acc_nl);
  assign nl_ln_1_if_251_acc_nl = conv_u2u_10_11(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:4])
      + 11'b11111111111;
  assign ln_1_if_251_acc_nl = nl_ln_1_if_251_acc_nl[10:0];
  assign ln_1_if_251_acc_itm_10_1 = readslicef_11_1_10(ln_1_if_251_acc_nl);
  assign nl_ln_1_if_250_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111111011;
  assign ln_1_if_250_acc_nl = nl_ln_1_if_250_acc_nl[12:0];
  assign ln_1_if_250_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_250_acc_nl);
  assign nl_ln_1_if_249_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:3])
      + 12'b111111111101;
  assign ln_1_if_249_acc_nl = nl_ln_1_if_249_acc_nl[11:0];
  assign ln_1_if_249_acc_itm_11_1 = readslicef_12_1_11(ln_1_if_249_acc_nl);
  assign nl_ln_1_if_248_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111111001;
  assign ln_1_if_248_acc_nl = nl_ln_1_if_248_acc_nl[12:0];
  assign ln_1_if_248_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_248_acc_nl);
  assign nl_ln_1_if_247_acc_nl = conv_u2u_9_10(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:5])
      + 10'b1111111111;
  assign ln_1_if_247_acc_nl = nl_ln_1_if_247_acc_nl[9:0];
  assign ln_1_if_247_acc_itm_9_1 = readslicef_10_1_9(ln_1_if_247_acc_nl);
  assign nl_ln_1_if_246_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111111011111;
  assign ln_1_if_246_acc_nl = nl_ln_1_if_246_acc_nl[14:0];
  assign ln_1_if_246_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_246_acc_nl);
  assign ln_1_nor_3_cse_1 = ~(ln_1_and_138_ssc_1 | ln_1_land_144_lpi_1_dfm_1);
  assign ln_1_nor_1_cse_1 = ~(ln_1_and_2_ssc_1 | ln_1_land_6_lpi_1_dfm_1);
  assign ln_1_land_8_lpi_1_dfm_1 = ln_1_if_7_acc_itm_5_1 & (~ ln_1_if_8_acc_itm_14_1);
  assign ln_1_land_9_lpi_1_dfm_1 = ln_1_if_8_acc_itm_14_1 & (~ ln_1_if_9_acc_itm_13_1);
  assign ln_1_land_11_lpi_1_dfm_1 = ln_1_if_10_acc_itm_14_1 & (~ ln_1_if_11_acc_itm_14_1);
  assign ln_1_land_13_lpi_1_dfm_1 = ln_1_if_12_acc_itm_10_1 & (~ ln_1_if_13_acc_itm_14_1);
  assign ln_1_land_15_lpi_1_dfm_1 = ln_1_if_14_acc_itm_13_1 & (~ ln_1_if_15_acc_itm_14_1);
  assign ln_1_and_4_ssc_1 = ln_1_if_6_acc_itm_8_1 & (~ ln_1_if_7_acc_itm_5_1) & (~(ln_1_land_9_lpi_1_dfm_1
      | ln_1_land_10_lpi_1_dfm_1)) & (~(ln_1_land_11_lpi_1_dfm_1 | ln_1_land_12_lpi_1_dfm_1))
      & (~(ln_1_land_13_lpi_1_dfm_1 | ln_1_land_14_lpi_1_dfm_1)) & (~(ln_1_land_15_lpi_1_dfm_1
      | ln_1_land_16_lpi_1_dfm_1)) & (~(ln_1_land_17_lpi_1_dfm_1 | ln_1_land_18_lpi_1_dfm_1))
      & (~(ln_1_land_19_lpi_1_dfm_1 | ln_1_land_20_lpi_1_dfm_1)) & (~(ln_1_land_21_lpi_1_dfm_1
      | ln_1_land_22_lpi_1_dfm_1)) & (~(ln_1_land_23_lpi_1_dfm_1 | ln_1_land_24_lpi_1_dfm_1))
      & (~(ln_1_land_25_lpi_1_dfm_1 | ln_1_land_26_lpi_1_dfm_1)) & (~(ln_1_land_27_lpi_1_dfm_1
      | ln_1_land_28_lpi_1_dfm_1)) & (~(ln_1_land_29_lpi_1_dfm_1 | ln_1_land_30_lpi_1_dfm_1))
      & (~(ln_1_land_31_lpi_1_dfm_1 | ln_1_land_32_lpi_1_dfm_1)) & (~(ln_1_land_33_lpi_1_dfm_1
      | ln_1_land_34_lpi_1_dfm_1)) & (~(ln_1_land_35_lpi_1_dfm_1 | ln_1_land_36_lpi_1_dfm_1))
      & (~(ln_1_land_37_lpi_1_dfm_1 | ln_1_land_38_lpi_1_dfm_1)) & (~(ln_1_land_39_lpi_1_dfm_1
      | ln_1_land_40_lpi_1_dfm_1)) & (~(ln_1_land_41_lpi_1_dfm_1 | ln_1_land_42_lpi_1_dfm_1))
      & (~(ln_1_land_43_lpi_1_dfm_1 | ln_1_land_44_lpi_1_dfm_1)) & (~(ln_1_land_45_lpi_1_dfm_1
      | ln_1_land_46_lpi_1_dfm_1)) & (~(ln_1_land_47_lpi_1_dfm_1 | ln_1_land_48_lpi_1_dfm_1
      | ln_1_land_49_lpi_1_dfm_1));
  assign ln_1_land_10_lpi_1_dfm_1 = ln_1_if_9_acc_itm_13_1 & (~ ln_1_if_10_acc_itm_14_1);
  assign ln_1_land_12_lpi_1_dfm_1 = ln_1_if_11_acc_itm_14_1 & (~ ln_1_if_12_acc_itm_10_1);
  assign ln_1_land_14_lpi_1_dfm_1 = ln_1_if_13_acc_itm_14_1 & (~ ln_1_if_14_acc_itm_13_1);
  assign ln_1_land_16_lpi_1_dfm_1 = ln_1_if_15_acc_itm_14_1 & (~ ln_1_if_16_acc_itm_12_1);
  assign ln_1_and_368_m1c_1 = (~(ln_1_land_229_lpi_1_dfm_1 | ln_1_land_230_lpi_1_dfm_1))
      & (~(ln_1_land_231_lpi_1_dfm_1 | ln_1_land_232_lpi_1_dfm_1)) & (~(ln_1_land_233_lpi_1_dfm_1
      | ln_1_land_234_lpi_1_dfm_1)) & (~(ln_1_land_235_lpi_1_dfm_1 | ln_1_land_236_lpi_1_dfm_1))
      & (~(ln_1_land_237_lpi_1_dfm_1 | ln_1_land_238_lpi_1_dfm_1)) & (~(ln_1_land_239_lpi_1_dfm_1
      | ln_1_land_240_lpi_1_dfm_1)) & (~(ln_1_land_241_lpi_1_dfm_1 | ln_1_land_242_lpi_1_dfm_1))
      & (~(ln_1_land_243_lpi_1_dfm_1 | ln_1_land_244_lpi_1_dfm_1));
  assign ln_1_land_4_lpi_1_dfm_1 = ln_1_if_3_acc_itm_6_1 & (~ ln_1_if_4_acc_itm_8_1);
  assign ln_1_and_2_ssc_1 = ln_1_if_4_acc_itm_8_1 & (~ ln_1_if_5_acc_itm_7_1);
  assign ln_1_land_6_lpi_1_dfm_1 = ln_1_if_5_acc_itm_7_1 & (~ ln_1_if_6_acc_itm_8_1);
  assign ln_1_nor_5_cse_1 = ~(ln_1_land_3_lpi_1_dfm_1 | ln_1_land_4_lpi_1_dfm_1);
  assign nl_ln_1_if_1_acc_nl = conv_u2u_7_8(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:7])
      + 8'b11111001;
  assign ln_1_if_1_acc_nl = nl_ln_1_if_1_acc_nl[7:0];
  assign ln_1_ret_13_0_lpi_1_dfm_257 = (readslicef_8_1_7(ln_1_if_1_acc_nl)) & (~
      ln_1_if_2_acc_itm_8_1);
  assign ln_1_land_3_lpi_1_dfm_1 = ln_1_if_2_acc_itm_8_1 & (~ ln_1_if_3_acc_itm_6_1);
  assign ln_1_ln_1_ln_1_nor_8_cse_1 = ~(ln_1_ret_13_0_lpi_1_dfm_257 | ln_1_land_4_lpi_1_dfm_1);
  assign nl_ln_1_if_144_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101111001;
  assign ln_1_if_144_acc_nl = nl_ln_1_if_144_acc_nl[14:0];
  assign ln_1_if_144_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_144_acc_nl);
  assign nl_ln_1_if_145_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111110111101;
  assign ln_1_if_145_acc_nl = nl_ln_1_if_145_acc_nl[13:0];
  assign ln_1_if_145_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_145_acc_nl);
  assign nl_ln_1_if_243_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111110111;
  assign ln_1_if_243_acc_nl = nl_ln_1_if_243_acc_nl[12:0];
  assign ln_1_if_243_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_243_acc_nl);
  assign nl_ln_1_if_242_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111111011011;
  assign ln_1_if_242_acc_nl = nl_ln_1_if_242_acc_nl[14:0];
  assign ln_1_if_242_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_242_acc_nl);
  assign nl_ln_1_if_241_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111101101;
  assign ln_1_if_241_acc_nl = nl_ln_1_if_241_acc_nl[13:0];
  assign ln_1_if_241_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_241_acc_nl);
  assign nl_ln_1_if_240_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111111011001;
  assign ln_1_if_240_acc_nl = nl_ln_1_if_240_acc_nl[14:0];
  assign ln_1_if_240_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_240_acc_nl);
  assign nl_ln_1_if_239_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:3])
      + 12'b111111111011;
  assign ln_1_if_239_acc_nl = nl_ln_1_if_239_acc_nl[11:0];
  assign ln_1_if_239_acc_itm_11_1 = readslicef_12_1_11(ln_1_if_239_acc_nl);
  assign nl_ln_1_if_238_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111111010111;
  assign ln_1_if_238_acc_nl = nl_ln_1_if_238_acc_nl[14:0];
  assign ln_1_if_238_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_238_acc_nl);
  assign nl_ln_1_if_237_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111101011;
  assign ln_1_if_237_acc_nl = nl_ln_1_if_237_acc_nl[13:0];
  assign ln_1_if_237_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_237_acc_nl);
  assign nl_ln_1_if_236_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111111010101;
  assign ln_1_if_236_acc_nl = nl_ln_1_if_236_acc_nl[14:0];
  assign ln_1_if_236_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_236_acc_nl);
  assign nl_ln_1_if_235_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111110101;
  assign ln_1_if_235_acc_nl = nl_ln_1_if_235_acc_nl[12:0];
  assign ln_1_if_235_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_235_acc_nl);
  assign nl_ln_1_if_234_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111111010011;
  assign ln_1_if_234_acc_nl = nl_ln_1_if_234_acc_nl[14:0];
  assign ln_1_if_234_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_234_acc_nl);
  assign nl_ln_1_if_233_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111101001;
  assign ln_1_if_233_acc_nl = nl_ln_1_if_233_acc_nl[13:0];
  assign ln_1_if_233_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_233_acc_nl);
  assign nl_ln_1_if_232_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111111010001;
  assign ln_1_if_232_acc_nl = nl_ln_1_if_232_acc_nl[14:0];
  assign ln_1_if_232_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_232_acc_nl);
  assign nl_ln_1_if_231_acc_nl = conv_u2u_10_11(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:4])
      + 11'b11111111101;
  assign ln_1_if_231_acc_nl = nl_ln_1_if_231_acc_nl[10:0];
  assign ln_1_if_231_acc_itm_10_1 = readslicef_11_1_10(ln_1_if_231_acc_nl);
  assign nl_ln_1_if_230_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111111001111;
  assign ln_1_if_230_acc_nl = nl_ln_1_if_230_acc_nl[14:0];
  assign ln_1_if_230_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_230_acc_nl);
  assign nl_ln_1_if_229_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111100111;
  assign ln_1_if_229_acc_nl = nl_ln_1_if_229_acc_nl[13:0];
  assign ln_1_if_229_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_229_acc_nl);
  assign nl_ln_1_if_228_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111111001101;
  assign ln_1_if_228_acc_nl = nl_ln_1_if_228_acc_nl[14:0];
  assign ln_1_if_228_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_228_acc_nl);
  assign nl_ln_1_if_227_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111110011;
  assign ln_1_if_227_acc_nl = nl_ln_1_if_227_acc_nl[12:0];
  assign ln_1_if_227_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_227_acc_nl);
  assign nl_ln_1_if_226_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111111001011;
  assign ln_1_if_226_acc_nl = nl_ln_1_if_226_acc_nl[14:0];
  assign ln_1_if_226_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_226_acc_nl);
  assign nl_ln_1_if_225_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111100101;
  assign ln_1_if_225_acc_nl = nl_ln_1_if_225_acc_nl[13:0];
  assign ln_1_if_225_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_225_acc_nl);
  assign nl_ln_1_if_224_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111111001001;
  assign ln_1_if_224_acc_nl = nl_ln_1_if_224_acc_nl[14:0];
  assign ln_1_if_224_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_224_acc_nl);
  assign nl_ln_1_if_223_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:3])
      + 12'b111111111001;
  assign ln_1_if_223_acc_nl = nl_ln_1_if_223_acc_nl[11:0];
  assign ln_1_if_223_acc_itm_11_1 = readslicef_12_1_11(ln_1_if_223_acc_nl);
  assign nl_ln_1_if_222_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111111000111;
  assign ln_1_if_222_acc_nl = nl_ln_1_if_222_acc_nl[14:0];
  assign ln_1_if_222_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_222_acc_nl);
  assign nl_ln_1_if_221_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111100011;
  assign ln_1_if_221_acc_nl = nl_ln_1_if_221_acc_nl[13:0];
  assign ln_1_if_221_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_221_acc_nl);
  assign nl_ln_1_if_220_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111111000101;
  assign ln_1_if_220_acc_nl = nl_ln_1_if_220_acc_nl[14:0];
  assign ln_1_if_220_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_220_acc_nl);
  assign nl_ln_1_if_219_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111110001;
  assign ln_1_if_219_acc_nl = nl_ln_1_if_219_acc_nl[12:0];
  assign ln_1_if_219_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_219_acc_nl);
  assign nl_ln_1_if_218_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111111000011;
  assign ln_1_if_218_acc_nl = nl_ln_1_if_218_acc_nl[14:0];
  assign ln_1_if_218_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_218_acc_nl);
  assign nl_ln_1_if_217_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111100001;
  assign ln_1_if_217_acc_nl = nl_ln_1_if_217_acc_nl[13:0];
  assign ln_1_if_217_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_217_acc_nl);
  assign nl_ln_1_if_216_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111111000001;
  assign ln_1_if_216_acc_nl = nl_ln_1_if_216_acc_nl[14:0];
  assign ln_1_if_216_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_216_acc_nl);
  assign nl_ln_1_if_215_acc_nl = conv_u2u_8_9(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:6])
      + 9'b111111111;
  assign ln_1_if_215_acc_nl = nl_ln_1_if_215_acc_nl[8:0];
  assign ln_1_if_215_acc_itm_8_1 = readslicef_9_1_8(ln_1_if_215_acc_nl);
  assign nl_ln_1_if_214_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110111111;
  assign ln_1_if_214_acc_nl = nl_ln_1_if_214_acc_nl[14:0];
  assign ln_1_if_214_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_214_acc_nl);
  assign nl_ln_1_if_213_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111011111;
  assign ln_1_if_213_acc_nl = nl_ln_1_if_213_acc_nl[13:0];
  assign ln_1_if_213_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_213_acc_nl);
  assign nl_ln_1_if_212_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110111101;
  assign ln_1_if_212_acc_nl = nl_ln_1_if_212_acc_nl[14:0];
  assign ln_1_if_212_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_212_acc_nl);
  assign nl_ln_1_if_211_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111101111;
  assign ln_1_if_211_acc_nl = nl_ln_1_if_211_acc_nl[12:0];
  assign ln_1_if_211_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_211_acc_nl);
  assign nl_ln_1_if_210_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110111011;
  assign ln_1_if_210_acc_nl = nl_ln_1_if_210_acc_nl[14:0];
  assign ln_1_if_210_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_210_acc_nl);
  assign nl_ln_1_if_209_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111011101;
  assign ln_1_if_209_acc_nl = nl_ln_1_if_209_acc_nl[13:0];
  assign ln_1_if_209_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_209_acc_nl);
  assign nl_ln_1_if_208_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110111001;
  assign ln_1_if_208_acc_nl = nl_ln_1_if_208_acc_nl[14:0];
  assign ln_1_if_208_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_208_acc_nl);
  assign nl_ln_1_if_207_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:3])
      + 12'b111111110111;
  assign ln_1_if_207_acc_nl = nl_ln_1_if_207_acc_nl[11:0];
  assign ln_1_if_207_acc_itm_11_1 = readslicef_12_1_11(ln_1_if_207_acc_nl);
  assign nl_ln_1_if_206_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110110111;
  assign ln_1_if_206_acc_nl = nl_ln_1_if_206_acc_nl[14:0];
  assign ln_1_if_206_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_206_acc_nl);
  assign nl_ln_1_if_205_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111011011;
  assign ln_1_if_205_acc_nl = nl_ln_1_if_205_acc_nl[13:0];
  assign ln_1_if_205_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_205_acc_nl);
  assign nl_ln_1_if_204_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110110101;
  assign ln_1_if_204_acc_nl = nl_ln_1_if_204_acc_nl[14:0];
  assign ln_1_if_204_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_204_acc_nl);
  assign nl_ln_1_if_203_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111101101;
  assign ln_1_if_203_acc_nl = nl_ln_1_if_203_acc_nl[12:0];
  assign ln_1_if_203_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_203_acc_nl);
  assign nl_ln_1_if_202_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110110011;
  assign ln_1_if_202_acc_nl = nl_ln_1_if_202_acc_nl[14:0];
  assign ln_1_if_202_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_202_acc_nl);
  assign nl_ln_1_if_201_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111011001;
  assign ln_1_if_201_acc_nl = nl_ln_1_if_201_acc_nl[13:0];
  assign ln_1_if_201_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_201_acc_nl);
  assign nl_ln_1_if_200_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110110001;
  assign ln_1_if_200_acc_nl = nl_ln_1_if_200_acc_nl[14:0];
  assign ln_1_if_200_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_200_acc_nl);
  assign nl_ln_1_if_199_acc_nl = conv_u2u_10_11(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:4])
      + 11'b11111111011;
  assign ln_1_if_199_acc_nl = nl_ln_1_if_199_acc_nl[10:0];
  assign ln_1_if_199_acc_itm_10_1 = readslicef_11_1_10(ln_1_if_199_acc_nl);
  assign nl_ln_1_if_198_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110101111;
  assign ln_1_if_198_acc_nl = nl_ln_1_if_198_acc_nl[14:0];
  assign ln_1_if_198_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_198_acc_nl);
  assign nl_ln_1_if_197_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111010111;
  assign ln_1_if_197_acc_nl = nl_ln_1_if_197_acc_nl[13:0];
  assign ln_1_if_197_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_197_acc_nl);
  assign nl_ln_1_if_196_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110101101;
  assign ln_1_if_196_acc_nl = nl_ln_1_if_196_acc_nl[14:0];
  assign ln_1_if_196_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_196_acc_nl);
  assign nl_ln_1_if_195_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111101011;
  assign ln_1_if_195_acc_nl = nl_ln_1_if_195_acc_nl[12:0];
  assign ln_1_if_195_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_195_acc_nl);
  assign nl_ln_1_if_194_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110101011;
  assign ln_1_if_194_acc_nl = nl_ln_1_if_194_acc_nl[14:0];
  assign ln_1_if_194_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_194_acc_nl);
  assign nl_ln_1_if_193_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111010101;
  assign ln_1_if_193_acc_nl = nl_ln_1_if_193_acc_nl[13:0];
  assign ln_1_if_193_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_193_acc_nl);
  assign nl_ln_1_if_192_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110101001;
  assign ln_1_if_192_acc_nl = nl_ln_1_if_192_acc_nl[14:0];
  assign ln_1_if_192_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_192_acc_nl);
  assign nl_ln_1_if_191_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:3])
      + 12'b111111110101;
  assign ln_1_if_191_acc_nl = nl_ln_1_if_191_acc_nl[11:0];
  assign ln_1_if_191_acc_itm_11_1 = readslicef_12_1_11(ln_1_if_191_acc_nl);
  assign nl_ln_1_if_190_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110100111;
  assign ln_1_if_190_acc_nl = nl_ln_1_if_190_acc_nl[14:0];
  assign ln_1_if_190_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_190_acc_nl);
  assign nl_ln_1_if_189_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111010011;
  assign ln_1_if_189_acc_nl = nl_ln_1_if_189_acc_nl[13:0];
  assign ln_1_if_189_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_189_acc_nl);
  assign nl_ln_1_if_188_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110100101;
  assign ln_1_if_188_acc_nl = nl_ln_1_if_188_acc_nl[14:0];
  assign ln_1_if_188_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_188_acc_nl);
  assign nl_ln_1_if_187_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111101001;
  assign ln_1_if_187_acc_nl = nl_ln_1_if_187_acc_nl[12:0];
  assign ln_1_if_187_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_187_acc_nl);
  assign nl_ln_1_if_186_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110100011;
  assign ln_1_if_186_acc_nl = nl_ln_1_if_186_acc_nl[14:0];
  assign ln_1_if_186_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_186_acc_nl);
  assign nl_ln_1_if_185_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111010001;
  assign ln_1_if_185_acc_nl = nl_ln_1_if_185_acc_nl[13:0];
  assign ln_1_if_185_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_185_acc_nl);
  assign nl_ln_1_if_184_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110100001;
  assign ln_1_if_184_acc_nl = nl_ln_1_if_184_acc_nl[14:0];
  assign ln_1_if_184_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_184_acc_nl);
  assign nl_ln_1_if_183_acc_nl = conv_u2u_9_10(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:5])
      + 10'b1111111101;
  assign ln_1_if_183_acc_nl = nl_ln_1_if_183_acc_nl[9:0];
  assign ln_1_if_183_acc_itm_9_1 = readslicef_10_1_9(ln_1_if_183_acc_nl);
  assign nl_ln_1_if_182_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110011111;
  assign ln_1_if_182_acc_nl = nl_ln_1_if_182_acc_nl[14:0];
  assign ln_1_if_182_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_182_acc_nl);
  assign nl_ln_1_if_181_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111001111;
  assign ln_1_if_181_acc_nl = nl_ln_1_if_181_acc_nl[13:0];
  assign ln_1_if_181_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_181_acc_nl);
  assign nl_ln_1_if_180_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110011101;
  assign ln_1_if_180_acc_nl = nl_ln_1_if_180_acc_nl[14:0];
  assign ln_1_if_180_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_180_acc_nl);
  assign nl_ln_1_if_179_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111100111;
  assign ln_1_if_179_acc_nl = nl_ln_1_if_179_acc_nl[12:0];
  assign ln_1_if_179_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_179_acc_nl);
  assign nl_ln_1_if_178_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110011011;
  assign ln_1_if_178_acc_nl = nl_ln_1_if_178_acc_nl[14:0];
  assign ln_1_if_178_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_178_acc_nl);
  assign nl_ln_1_if_177_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111001101;
  assign ln_1_if_177_acc_nl = nl_ln_1_if_177_acc_nl[13:0];
  assign ln_1_if_177_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_177_acc_nl);
  assign nl_ln_1_if_176_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110011001;
  assign ln_1_if_176_acc_nl = nl_ln_1_if_176_acc_nl[14:0];
  assign ln_1_if_176_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_176_acc_nl);
  assign nl_ln_1_if_175_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:3])
      + 12'b111111110011;
  assign ln_1_if_175_acc_nl = nl_ln_1_if_175_acc_nl[11:0];
  assign ln_1_if_175_acc_itm_11_1 = readslicef_12_1_11(ln_1_if_175_acc_nl);
  assign nl_ln_1_if_174_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110010111;
  assign ln_1_if_174_acc_nl = nl_ln_1_if_174_acc_nl[14:0];
  assign ln_1_if_174_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_174_acc_nl);
  assign nl_ln_1_if_173_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111001011;
  assign ln_1_if_173_acc_nl = nl_ln_1_if_173_acc_nl[13:0];
  assign ln_1_if_173_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_173_acc_nl);
  assign nl_ln_1_if_172_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110010101;
  assign ln_1_if_172_acc_nl = nl_ln_1_if_172_acc_nl[14:0];
  assign ln_1_if_172_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_172_acc_nl);
  assign nl_ln_1_if_171_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111100101;
  assign ln_1_if_171_acc_nl = nl_ln_1_if_171_acc_nl[12:0];
  assign ln_1_if_171_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_171_acc_nl);
  assign nl_ln_1_if_170_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110010011;
  assign ln_1_if_170_acc_nl = nl_ln_1_if_170_acc_nl[14:0];
  assign ln_1_if_170_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_170_acc_nl);
  assign nl_ln_1_if_169_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111001001;
  assign ln_1_if_169_acc_nl = nl_ln_1_if_169_acc_nl[13:0];
  assign ln_1_if_169_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_169_acc_nl);
  assign nl_ln_1_if_168_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110010001;
  assign ln_1_if_168_acc_nl = nl_ln_1_if_168_acc_nl[14:0];
  assign ln_1_if_168_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_168_acc_nl);
  assign nl_ln_1_if_167_acc_nl = conv_u2u_10_11(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:4])
      + 11'b11111111001;
  assign ln_1_if_167_acc_nl = nl_ln_1_if_167_acc_nl[10:0];
  assign ln_1_if_167_acc_itm_10_1 = readslicef_11_1_10(ln_1_if_167_acc_nl);
  assign nl_ln_1_if_166_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110001111;
  assign ln_1_if_166_acc_nl = nl_ln_1_if_166_acc_nl[14:0];
  assign ln_1_if_166_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_166_acc_nl);
  assign nl_ln_1_if_165_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111000111;
  assign ln_1_if_165_acc_nl = nl_ln_1_if_165_acc_nl[13:0];
  assign ln_1_if_165_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_165_acc_nl);
  assign nl_ln_1_if_164_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110001101;
  assign ln_1_if_164_acc_nl = nl_ln_1_if_164_acc_nl[14:0];
  assign ln_1_if_164_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_164_acc_nl);
  assign nl_ln_1_if_163_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111100011;
  assign ln_1_if_163_acc_nl = nl_ln_1_if_163_acc_nl[12:0];
  assign ln_1_if_163_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_163_acc_nl);
  assign nl_ln_1_if_162_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110001011;
  assign ln_1_if_162_acc_nl = nl_ln_1_if_162_acc_nl[14:0];
  assign ln_1_if_162_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_162_acc_nl);
  assign nl_ln_1_if_161_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111000101;
  assign ln_1_if_161_acc_nl = nl_ln_1_if_161_acc_nl[13:0];
  assign ln_1_if_161_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_161_acc_nl);
  assign nl_ln_1_if_160_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110001001;
  assign ln_1_if_160_acc_nl = nl_ln_1_if_160_acc_nl[14:0];
  assign ln_1_if_160_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_160_acc_nl);
  assign nl_ln_1_if_159_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:3])
      + 12'b111111110001;
  assign ln_1_if_159_acc_nl = nl_ln_1_if_159_acc_nl[11:0];
  assign ln_1_if_159_acc_itm_11_1 = readslicef_12_1_11(ln_1_if_159_acc_nl);
  assign nl_ln_1_if_158_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110000111;
  assign ln_1_if_158_acc_nl = nl_ln_1_if_158_acc_nl[14:0];
  assign ln_1_if_158_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_158_acc_nl);
  assign nl_ln_1_if_157_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111000011;
  assign ln_1_if_157_acc_nl = nl_ln_1_if_157_acc_nl[13:0];
  assign ln_1_if_157_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_157_acc_nl);
  assign nl_ln_1_if_156_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110000101;
  assign ln_1_if_156_acc_nl = nl_ln_1_if_156_acc_nl[14:0];
  assign ln_1_if_156_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_156_acc_nl);
  assign nl_ln_1_if_155_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111100001;
  assign ln_1_if_155_acc_nl = nl_ln_1_if_155_acc_nl[12:0];
  assign ln_1_if_155_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_155_acc_nl);
  assign nl_ln_1_if_154_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110000011;
  assign ln_1_if_154_acc_nl = nl_ln_1_if_154_acc_nl[14:0];
  assign ln_1_if_154_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_154_acc_nl);
  assign nl_ln_1_if_153_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111111000001;
  assign ln_1_if_153_acc_nl = nl_ln_1_if_153_acc_nl[13:0];
  assign ln_1_if_153_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_153_acc_nl);
  assign nl_ln_1_if_152_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111110000001;
  assign ln_1_if_152_acc_nl = nl_ln_1_if_152_acc_nl[14:0];
  assign ln_1_if_152_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_152_acc_nl);
  assign nl_ln_1_if_151_acc_nl = conv_u2u_7_8(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:7])
      + 8'b11111111;
  assign ln_1_if_151_acc_nl = nl_ln_1_if_151_acc_nl[7:0];
  assign ln_1_if_151_acc_itm_7_1 = readslicef_8_1_7(ln_1_if_151_acc_nl);
  assign nl_ln_1_if_150_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101111111;
  assign ln_1_if_150_acc_nl = nl_ln_1_if_150_acc_nl[14:0];
  assign ln_1_if_150_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_150_acc_nl);
  assign nl_ln_1_if_149_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111110111111;
  assign ln_1_if_149_acc_nl = nl_ln_1_if_149_acc_nl[13:0];
  assign ln_1_if_149_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_149_acc_nl);
  assign nl_ln_1_if_148_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101111101;
  assign ln_1_if_148_acc_nl = nl_ln_1_if_148_acc_nl[14:0];
  assign ln_1_if_148_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_148_acc_nl);
  assign nl_ln_1_if_147_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111011111;
  assign ln_1_if_147_acc_nl = nl_ln_1_if_147_acc_nl[12:0];
  assign ln_1_if_147_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_147_acc_nl);
  assign nl_ln_1_if_146_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101111011;
  assign ln_1_if_146_acc_nl = nl_ln_1_if_146_acc_nl[14:0];
  assign ln_1_if_146_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_146_acc_nl);
  assign nl_ln_1_if_142_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101110111;
  assign ln_1_if_142_acc_nl = nl_ln_1_if_142_acc_nl[14:0];
  assign ln_1_if_142_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_142_acc_nl);
  assign nl_ln_1_if_143_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:3])
      + 12'b111111101111;
  assign ln_1_if_143_acc_nl = nl_ln_1_if_143_acc_nl[11:0];
  assign ln_1_if_143_acc_itm_11_1 = readslicef_12_1_11(ln_1_if_143_acc_nl);
  assign nl_ln_1_if_141_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111110111011;
  assign ln_1_if_141_acc_nl = nl_ln_1_if_141_acc_nl[13:0];
  assign ln_1_if_141_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_141_acc_nl);
  assign nl_ln_1_if_140_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101110101;
  assign ln_1_if_140_acc_nl = nl_ln_1_if_140_acc_nl[14:0];
  assign ln_1_if_140_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_140_acc_nl);
  assign nl_ln_1_if_52_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111010001101;
  assign ln_1_if_52_acc_nl = nl_ln_1_if_52_acc_nl[14:0];
  assign ln_1_if_52_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_52_acc_nl);
  assign nl_ln_1_if_53_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111010010001;
  assign ln_1_if_53_acc_nl = nl_ln_1_if_53_acc_nl[14:0];
  assign ln_1_if_53_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_53_acc_nl);
  assign nl_ln_1_if_49_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111110100001;
  assign ln_1_if_49_acc_nl = nl_ln_1_if_49_acc_nl[12:0];
  assign ln_1_if_49_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_49_acc_nl);
  assign nl_ln_1_if_50_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111010000111;
  assign ln_1_if_50_acc_nl = nl_ln_1_if_50_acc_nl[14:0];
  assign ln_1_if_50_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_50_acc_nl);
  assign nl_ln_1_if_6_acc_nl = conv_u2u_8_9(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:6])
      + 9'b111110111;
  assign ln_1_if_6_acc_nl = nl_ln_1_if_6_acc_nl[8:0];
  assign ln_1_if_6_acc_itm_8_1 = readslicef_9_1_8(ln_1_if_6_acc_nl);
  assign nl_ln_1_if_7_acc_nl = conv_u2u_5_6(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:9])
      + 6'b111111;
  assign ln_1_if_7_acc_nl = nl_ln_1_if_7_acc_nl[5:0];
  assign ln_1_if_7_acc_itm_5_1 = readslicef_6_1_5(ln_1_if_7_acc_nl);
  assign nl_ln_1_if_139_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111011101;
  assign ln_1_if_139_acc_nl = nl_ln_1_if_139_acc_nl[12:0];
  assign ln_1_if_139_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_139_acc_nl);
  assign nl_ln_1_if_138_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101110011;
  assign ln_1_if_138_acc_nl = nl_ln_1_if_138_acc_nl[14:0];
  assign ln_1_if_138_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_138_acc_nl);
  assign nl_ln_1_if_137_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111110111001;
  assign ln_1_if_137_acc_nl = nl_ln_1_if_137_acc_nl[13:0];
  assign ln_1_if_137_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_137_acc_nl);
  assign nl_ln_1_if_136_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101110001;
  assign ln_1_if_136_acc_nl = nl_ln_1_if_136_acc_nl[14:0];
  assign ln_1_if_136_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_136_acc_nl);
  assign nl_ln_1_if_135_acc_nl = conv_u2u_10_11(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:4])
      + 11'b11111110111;
  assign ln_1_if_135_acc_nl = nl_ln_1_if_135_acc_nl[10:0];
  assign ln_1_if_135_acc_itm_10_1 = readslicef_11_1_10(ln_1_if_135_acc_nl);
  assign nl_ln_1_if_134_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101101111;
  assign ln_1_if_134_acc_nl = nl_ln_1_if_134_acc_nl[14:0];
  assign ln_1_if_134_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_134_acc_nl);
  assign nl_ln_1_if_133_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111110110111;
  assign ln_1_if_133_acc_nl = nl_ln_1_if_133_acc_nl[13:0];
  assign ln_1_if_133_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_133_acc_nl);
  assign nl_ln_1_if_132_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101101101;
  assign ln_1_if_132_acc_nl = nl_ln_1_if_132_acc_nl[14:0];
  assign ln_1_if_132_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_132_acc_nl);
  assign nl_ln_1_if_131_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111011011;
  assign ln_1_if_131_acc_nl = nl_ln_1_if_131_acc_nl[12:0];
  assign ln_1_if_131_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_131_acc_nl);
  assign nl_ln_1_if_130_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101101011;
  assign ln_1_if_130_acc_nl = nl_ln_1_if_130_acc_nl[14:0];
  assign ln_1_if_130_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_130_acc_nl);
  assign nl_ln_1_if_129_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111110110101;
  assign ln_1_if_129_acc_nl = nl_ln_1_if_129_acc_nl[13:0];
  assign ln_1_if_129_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_129_acc_nl);
  assign nl_ln_1_if_128_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101101001;
  assign ln_1_if_128_acc_nl = nl_ln_1_if_128_acc_nl[14:0];
  assign ln_1_if_128_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_128_acc_nl);
  assign nl_ln_1_if_127_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:3])
      + 12'b111111101101;
  assign ln_1_if_127_acc_nl = nl_ln_1_if_127_acc_nl[11:0];
  assign ln_1_if_127_acc_itm_11_1 = readslicef_12_1_11(ln_1_if_127_acc_nl);
  assign nl_ln_1_if_126_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101100111;
  assign ln_1_if_126_acc_nl = nl_ln_1_if_126_acc_nl[14:0];
  assign ln_1_if_126_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_126_acc_nl);
  assign nl_ln_1_if_125_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111110110011;
  assign ln_1_if_125_acc_nl = nl_ln_1_if_125_acc_nl[13:0];
  assign ln_1_if_125_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_125_acc_nl);
  assign nl_ln_1_if_124_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101100101;
  assign ln_1_if_124_acc_nl = nl_ln_1_if_124_acc_nl[14:0];
  assign ln_1_if_124_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_124_acc_nl);
  assign nl_ln_1_if_123_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111011001;
  assign ln_1_if_123_acc_nl = nl_ln_1_if_123_acc_nl[12:0];
  assign ln_1_if_123_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_123_acc_nl);
  assign nl_ln_1_if_122_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101100011;
  assign ln_1_if_122_acc_nl = nl_ln_1_if_122_acc_nl[14:0];
  assign ln_1_if_122_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_122_acc_nl);
  assign nl_ln_1_if_121_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111110110001;
  assign ln_1_if_121_acc_nl = nl_ln_1_if_121_acc_nl[13:0];
  assign ln_1_if_121_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_121_acc_nl);
  assign nl_ln_1_if_120_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101100001;
  assign ln_1_if_120_acc_nl = nl_ln_1_if_120_acc_nl[14:0];
  assign ln_1_if_120_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_120_acc_nl);
  assign nl_ln_1_if_119_acc_nl = conv_u2u_9_10(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:5])
      + 10'b1111111011;
  assign ln_1_if_119_acc_nl = nl_ln_1_if_119_acc_nl[9:0];
  assign ln_1_if_119_acc_itm_9_1 = readslicef_10_1_9(ln_1_if_119_acc_nl);
  assign nl_ln_1_if_118_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101011101;
  assign ln_1_if_118_acc_nl = nl_ln_1_if_118_acc_nl[14:0];
  assign ln_1_if_118_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_118_acc_nl);
  assign nl_ln_1_if_117_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111110101101;
  assign ln_1_if_117_acc_nl = nl_ln_1_if_117_acc_nl[13:0];
  assign ln_1_if_117_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_117_acc_nl);
  assign nl_ln_1_if_116_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101010111;
  assign ln_1_if_116_acc_nl = nl_ln_1_if_116_acc_nl[14:0];
  assign ln_1_if_116_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_116_acc_nl);
  assign nl_ln_1_if_115_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101010011;
  assign ln_1_if_115_acc_nl = nl_ln_1_if_115_acc_nl[14:0];
  assign ln_1_if_115_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_115_acc_nl);
  assign nl_ln_1_if_114_acc_nl = conv_u2u_10_11(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:4])
      + 11'b11111110101;
  assign ln_1_if_114_acc_nl = nl_ln_1_if_114_acc_nl[10:0];
  assign ln_1_if_114_acc_itm_10_1 = readslicef_11_1_10(ln_1_if_114_acc_nl);
  assign nl_ln_1_if_113_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101001101;
  assign ln_1_if_113_acc_nl = nl_ln_1_if_113_acc_nl[14:0];
  assign ln_1_if_113_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_113_acc_nl);
  assign nl_ln_1_if_112_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111110100101;
  assign ln_1_if_112_acc_nl = nl_ln_1_if_112_acc_nl[13:0];
  assign ln_1_if_112_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_112_acc_nl);
  assign nl_ln_1_if_111_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101000111;
  assign ln_1_if_111_acc_nl = nl_ln_1_if_111_acc_nl[14:0];
  assign ln_1_if_111_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_111_acc_nl);
  assign nl_ln_1_if_110_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111010001;
  assign ln_1_if_110_acc_nl = nl_ln_1_if_110_acc_nl[12:0];
  assign ln_1_if_110_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_110_acc_nl);
  assign nl_ln_1_if_109_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111101000001;
  assign ln_1_if_109_acc_nl = nl_ln_1_if_109_acc_nl[14:0];
  assign ln_1_if_109_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_109_acc_nl);
  assign nl_ln_1_if_108_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111100111101;
  assign ln_1_if_108_acc_nl = nl_ln_1_if_108_acc_nl[14:0];
  assign ln_1_if_108_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_108_acc_nl);
  assign nl_ln_1_if_107_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111110011101;
  assign ln_1_if_107_acc_nl = nl_ln_1_if_107_acc_nl[13:0];
  assign ln_1_if_107_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_107_acc_nl);
  assign nl_ln_1_if_106_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111100110111;
  assign ln_1_if_106_acc_nl = nl_ln_1_if_106_acc_nl[14:0];
  assign ln_1_if_106_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_106_acc_nl);
  assign nl_ln_1_if_105_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111001101;
  assign ln_1_if_105_acc_nl = nl_ln_1_if_105_acc_nl[12:0];
  assign ln_1_if_105_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_105_acc_nl);
  assign nl_ln_1_if_104_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111100110001;
  assign ln_1_if_104_acc_nl = nl_ln_1_if_104_acc_nl[14:0];
  assign ln_1_if_104_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_104_acc_nl);
  assign nl_ln_1_if_103_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111110010111;
  assign ln_1_if_103_acc_nl = nl_ln_1_if_103_acc_nl[13:0];
  assign ln_1_if_103_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_103_acc_nl);
  assign nl_ln_1_if_102_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111100101011;
  assign ln_1_if_102_acc_nl = nl_ln_1_if_102_acc_nl[14:0];
  assign ln_1_if_102_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_102_acc_nl);
  assign nl_ln_1_if_101_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111100100111;
  assign ln_1_if_101_acc_nl = nl_ln_1_if_101_acc_nl[14:0];
  assign ln_1_if_101_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_101_acc_nl);
  assign nl_ln_1_if_100_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111111001001;
  assign ln_1_if_100_acc_nl = nl_ln_1_if_100_acc_nl[12:0];
  assign ln_1_if_100_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_100_acc_nl);
  assign nl_ln_1_if_99_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111100100001;
  assign ln_1_if_99_acc_nl = nl_ln_1_if_99_acc_nl[14:0];
  assign ln_1_if_99_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_99_acc_nl);
  assign nl_ln_1_if_98_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111110001111;
  assign ln_1_if_98_acc_nl = nl_ln_1_if_98_acc_nl[13:0];
  assign ln_1_if_98_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_98_acc_nl);
  assign nl_ln_1_if_97_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111100011011;
  assign ln_1_if_97_acc_nl = nl_ln_1_if_97_acc_nl[14:0];
  assign ln_1_if_97_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_97_acc_nl);
  assign nl_ln_1_if_96_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:3])
      + 12'b111111100011;
  assign ln_1_if_96_acc_nl = nl_ln_1_if_96_acc_nl[11:0];
  assign ln_1_if_96_acc_itm_11_1 = readslicef_12_1_11(ln_1_if_96_acc_nl);
  assign nl_ln_1_if_95_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111100010101;
  assign ln_1_if_95_acc_nl = nl_ln_1_if_95_acc_nl[14:0];
  assign ln_1_if_95_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_95_acc_nl);
  assign nl_ln_1_if_94_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111100010001;
  assign ln_1_if_94_acc_nl = nl_ln_1_if_94_acc_nl[14:0];
  assign ln_1_if_94_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_94_acc_nl);
  assign nl_ln_1_if_93_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111110000111;
  assign ln_1_if_93_acc_nl = nl_ln_1_if_93_acc_nl[13:0];
  assign ln_1_if_93_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_93_acc_nl);
  assign nl_ln_1_if_92_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111100001011;
  assign ln_1_if_92_acc_nl = nl_ln_1_if_92_acc_nl[14:0];
  assign ln_1_if_92_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_92_acc_nl);
  assign nl_ln_1_if_91_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:3])
      + 12'b111111100001;
  assign ln_1_if_91_acc_nl = nl_ln_1_if_91_acc_nl[11:0];
  assign ln_1_if_91_acc_itm_11_1 = readslicef_12_1_11(ln_1_if_91_acc_nl);
  assign nl_ln_1_if_90_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111100000101;
  assign ln_1_if_90_acc_nl = nl_ln_1_if_90_acc_nl[14:0];
  assign ln_1_if_90_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_90_acc_nl);
  assign nl_ln_1_if_89_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111110000001;
  assign ln_1_if_89_acc_nl = nl_ln_1_if_89_acc_nl[13:0];
  assign ln_1_if_89_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_89_acc_nl);
  assign nl_ln_1_if_88_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111011111111;
  assign ln_1_if_88_acc_nl = nl_ln_1_if_88_acc_nl[14:0];
  assign ln_1_if_88_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_88_acc_nl);
  assign nl_ln_1_if_87_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111011111011;
  assign ln_1_if_87_acc_nl = nl_ln_1_if_87_acc_nl[14:0];
  assign ln_1_if_87_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_87_acc_nl);
  assign nl_ln_1_if_86_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:3])
      + 12'b111111011111;
  assign ln_1_if_86_acc_nl = nl_ln_1_if_86_acc_nl[11:0];
  assign ln_1_if_86_acc_itm_11_1 = readslicef_12_1_11(ln_1_if_86_acc_nl);
  assign nl_ln_1_if_85_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111011110101;
  assign ln_1_if_85_acc_nl = nl_ln_1_if_85_acc_nl[14:0];
  assign ln_1_if_85_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_85_acc_nl);
  assign nl_ln_1_if_84_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111101111001;
  assign ln_1_if_84_acc_nl = nl_ln_1_if_84_acc_nl[13:0];
  assign ln_1_if_84_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_84_acc_nl);
  assign nl_ln_1_if_83_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111011101111;
  assign ln_1_if_83_acc_nl = nl_ln_1_if_83_acc_nl[14:0];
  assign ln_1_if_83_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_83_acc_nl);
  assign nl_ln_1_if_82_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111110111011;
  assign ln_1_if_82_acc_nl = nl_ln_1_if_82_acc_nl[12:0];
  assign ln_1_if_82_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_82_acc_nl);
  assign nl_ln_1_if_81_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111011101001;
  assign ln_1_if_81_acc_nl = nl_ln_1_if_81_acc_nl[14:0];
  assign ln_1_if_81_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_81_acc_nl);
  assign nl_ln_1_if_80_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111011100101;
  assign ln_1_if_80_acc_nl = nl_ln_1_if_80_acc_nl[14:0];
  assign ln_1_if_80_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_80_acc_nl);
  assign nl_ln_1_if_79_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111101110001;
  assign ln_1_if_79_acc_nl = nl_ln_1_if_79_acc_nl[13:0];
  assign ln_1_if_79_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_79_acc_nl);
  assign nl_ln_1_if_78_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111011011111;
  assign ln_1_if_78_acc_nl = nl_ln_1_if_78_acc_nl[14:0];
  assign ln_1_if_78_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_78_acc_nl);
  assign nl_ln_1_if_77_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111110110111;
  assign ln_1_if_77_acc_nl = nl_ln_1_if_77_acc_nl[12:0];
  assign ln_1_if_77_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_77_acc_nl);
  assign nl_ln_1_if_76_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111011011001;
  assign ln_1_if_76_acc_nl = nl_ln_1_if_76_acc_nl[14:0];
  assign ln_1_if_76_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_76_acc_nl);
  assign nl_ln_1_if_75_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111101101011;
  assign ln_1_if_75_acc_nl = nl_ln_1_if_75_acc_nl[13:0];
  assign ln_1_if_75_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_75_acc_nl);
  assign nl_ln_1_if_74_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111011010011;
  assign ln_1_if_74_acc_nl = nl_ln_1_if_74_acc_nl[14:0];
  assign ln_1_if_74_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_74_acc_nl);
  assign nl_ln_1_if_73_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111011001111;
  assign ln_1_if_73_acc_nl = nl_ln_1_if_73_acc_nl[14:0];
  assign ln_1_if_73_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_73_acc_nl);
  assign nl_ln_1_if_72_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111110110011;
  assign ln_1_if_72_acc_nl = nl_ln_1_if_72_acc_nl[12:0];
  assign ln_1_if_72_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_72_acc_nl);
  assign nl_ln_1_if_71_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111011001001;
  assign ln_1_if_71_acc_nl = nl_ln_1_if_71_acc_nl[14:0];
  assign ln_1_if_71_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_71_acc_nl);
  assign nl_ln_1_if_70_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111101100011;
  assign ln_1_if_70_acc_nl = nl_ln_1_if_70_acc_nl[13:0];
  assign ln_1_if_70_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_70_acc_nl);
  assign nl_ln_1_if_69_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111011000011;
  assign ln_1_if_69_acc_nl = nl_ln_1_if_69_acc_nl[14:0];
  assign ln_1_if_69_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_69_acc_nl);
  assign nl_ln_1_if_68_acc_nl = conv_u2u_8_9(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:6])
      + 9'b111111011;
  assign ln_1_if_68_acc_nl = nl_ln_1_if_68_acc_nl[8:0];
  assign ln_1_if_68_acc_itm_8_1 = readslicef_9_1_8(ln_1_if_68_acc_nl);
  assign nl_ln_1_if_67_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111010111101;
  assign ln_1_if_67_acc_nl = nl_ln_1_if_67_acc_nl[14:0];
  assign ln_1_if_67_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_67_acc_nl);
  assign nl_ln_1_if_66_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111010111001;
  assign ln_1_if_66_acc_nl = nl_ln_1_if_66_acc_nl[14:0];
  assign ln_1_if_66_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_66_acc_nl);
  assign nl_ln_1_if_65_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111101011011;
  assign ln_1_if_65_acc_nl = nl_ln_1_if_65_acc_nl[13:0];
  assign ln_1_if_65_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_65_acc_nl);
  assign nl_ln_1_if_64_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111010110011;
  assign ln_1_if_64_acc_nl = nl_ln_1_if_64_acc_nl[14:0];
  assign ln_1_if_64_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_64_acc_nl);
  assign nl_ln_1_if_63_acc_nl = conv_u2u_10_11(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:4])
      + 11'b11111101011;
  assign ln_1_if_63_acc_nl = nl_ln_1_if_63_acc_nl[10:0];
  assign ln_1_if_63_acc_itm_10_1 = readslicef_11_1_10(ln_1_if_63_acc_nl);
  assign nl_ln_1_if_62_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111010101101;
  assign ln_1_if_62_acc_nl = nl_ln_1_if_62_acc_nl[14:0];
  assign ln_1_if_62_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_62_acc_nl);
  assign nl_ln_1_if_61_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111101010101;
  assign ln_1_if_61_acc_nl = nl_ln_1_if_61_acc_nl[13:0];
  assign ln_1_if_61_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_61_acc_nl);
  assign nl_ln_1_if_60_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111010100111;
  assign ln_1_if_60_acc_nl = nl_ln_1_if_60_acc_nl[14:0];
  assign ln_1_if_60_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_60_acc_nl);
  assign nl_ln_1_if_59_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111010100011;
  assign ln_1_if_59_acc_nl = nl_ln_1_if_59_acc_nl[14:0];
  assign ln_1_if_59_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_59_acc_nl);
  assign nl_ln_1_if_58_acc_nl = conv_u2u_9_10(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:5])
      + 10'b1111110101;
  assign ln_1_if_58_acc_nl = nl_ln_1_if_58_acc_nl[9:0];
  assign ln_1_if_58_acc_itm_9_1 = readslicef_10_1_9(ln_1_if_58_acc_nl);
  assign nl_ln_1_if_57_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111010011101;
  assign ln_1_if_57_acc_nl = nl_ln_1_if_57_acc_nl[14:0];
  assign ln_1_if_57_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_57_acc_nl);
  assign nl_ln_1_if_56_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111101001101;
  assign ln_1_if_56_acc_nl = nl_ln_1_if_56_acc_nl[13:0];
  assign ln_1_if_56_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_56_acc_nl);
  assign nl_ln_1_if_55_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111010010111;
  assign ln_1_if_55_acc_nl = nl_ln_1_if_55_acc_nl[14:0];
  assign ln_1_if_55_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_55_acc_nl);
  assign nl_ln_1_if_54_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111110100101;
  assign ln_1_if_54_acc_nl = nl_ln_1_if_54_acc_nl[12:0];
  assign ln_1_if_54_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_54_acc_nl);
  assign nl_ln_1_if_51_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111101000101;
  assign ln_1_if_51_acc_nl = nl_ln_1_if_51_acc_nl[13:0];
  assign ln_1_if_51_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_51_acc_nl);
  assign nl_ln_1_if_48_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111010000001;
  assign ln_1_if_48_acc_nl = nl_ln_1_if_48_acc_nl[14:0];
  assign ln_1_if_48_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_48_acc_nl);
  assign nl_ln_1_if_47_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111100111111;
  assign ln_1_if_47_acc_nl = nl_ln_1_if_47_acc_nl[13:0];
  assign ln_1_if_47_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_47_acc_nl);
  assign nl_ln_1_if_46_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111001111011;
  assign ln_1_if_46_acc_nl = nl_ln_1_if_46_acc_nl[14:0];
  assign ln_1_if_46_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_46_acc_nl);
  assign nl_ln_1_if_45_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111001110111;
  assign ln_1_if_45_acc_nl = nl_ln_1_if_45_acc_nl[14:0];
  assign ln_1_if_45_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_45_acc_nl);
  assign nl_ln_1_if_44_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111110011101;
  assign ln_1_if_44_acc_nl = nl_ln_1_if_44_acc_nl[12:0];
  assign ln_1_if_44_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_44_acc_nl);
  assign nl_ln_1_if_43_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111001110001;
  assign ln_1_if_43_acc_nl = nl_ln_1_if_43_acc_nl[14:0];
  assign ln_1_if_43_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_43_acc_nl);
  assign nl_ln_1_if_42_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111100110111;
  assign ln_1_if_42_acc_nl = nl_ln_1_if_42_acc_nl[13:0];
  assign ln_1_if_42_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_42_acc_nl);
  assign nl_ln_1_if_41_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111001101011;
  assign ln_1_if_41_acc_nl = nl_ln_1_if_41_acc_nl[14:0];
  assign ln_1_if_41_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_41_acc_nl);
  assign nl_ln_1_if_40_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:3])
      + 12'b111111001101;
  assign ln_1_if_40_acc_nl = nl_ln_1_if_40_acc_nl[11:0];
  assign ln_1_if_40_acc_itm_11_1 = readslicef_12_1_11(ln_1_if_40_acc_nl);
  assign nl_ln_1_if_39_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111001100101;
  assign ln_1_if_39_acc_nl = nl_ln_1_if_39_acc_nl[14:0];
  assign ln_1_if_39_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_39_acc_nl);
  assign nl_ln_1_if_38_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111001100001;
  assign ln_1_if_38_acc_nl = nl_ln_1_if_38_acc_nl[14:0];
  assign ln_1_if_38_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_38_acc_nl);
  assign nl_ln_1_if_37_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111100101111;
  assign ln_1_if_37_acc_nl = nl_ln_1_if_37_acc_nl[13:0];
  assign ln_1_if_37_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_37_acc_nl);
  assign nl_ln_1_if_36_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111001011011;
  assign ln_1_if_36_acc_nl = nl_ln_1_if_36_acc_nl[14:0];
  assign ln_1_if_36_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_36_acc_nl);
  assign nl_ln_1_if_35_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:3])
      + 12'b111111001011;
  assign ln_1_if_35_acc_nl = nl_ln_1_if_35_acc_nl[11:0];
  assign ln_1_if_35_acc_itm_11_1 = readslicef_12_1_11(ln_1_if_35_acc_nl);
  assign nl_ln_1_if_34_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111001010101;
  assign ln_1_if_34_acc_nl = nl_ln_1_if_34_acc_nl[14:0];
  assign ln_1_if_34_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_34_acc_nl);
  assign nl_ln_1_if_33_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111100101001;
  assign ln_1_if_33_acc_nl = nl_ln_1_if_33_acc_nl[13:0];
  assign ln_1_if_33_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_33_acc_nl);
  assign nl_ln_1_if_32_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111001001111;
  assign ln_1_if_32_acc_nl = nl_ln_1_if_32_acc_nl[14:0];
  assign ln_1_if_32_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_32_acc_nl);
  assign nl_ln_1_if_31_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111001001011;
  assign ln_1_if_31_acc_nl = nl_ln_1_if_31_acc_nl[14:0];
  assign ln_1_if_31_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_31_acc_nl);
  assign nl_ln_1_if_30_acc_nl = conv_u2u_11_12(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:3])
      + 12'b111111001001;
  assign ln_1_if_30_acc_nl = nl_ln_1_if_30_acc_nl[11:0];
  assign ln_1_if_30_acc_itm_11_1 = readslicef_12_1_11(ln_1_if_30_acc_nl);
  assign nl_ln_1_if_29_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111001000101;
  assign ln_1_if_29_acc_nl = nl_ln_1_if_29_acc_nl[14:0];
  assign ln_1_if_29_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_29_acc_nl);
  assign nl_ln_1_if_28_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111100100001;
  assign ln_1_if_28_acc_nl = nl_ln_1_if_28_acc_nl[13:0];
  assign ln_1_if_28_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_28_acc_nl);
  assign nl_ln_1_if_27_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111000111111;
  assign ln_1_if_27_acc_nl = nl_ln_1_if_27_acc_nl[14:0];
  assign ln_1_if_27_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_27_acc_nl);
  assign nl_ln_1_if_26_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111110001111;
  assign ln_1_if_26_acc_nl = nl_ln_1_if_26_acc_nl[12:0];
  assign ln_1_if_26_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_26_acc_nl);
  assign nl_ln_1_if_25_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111000111001;
  assign ln_1_if_25_acc_nl = nl_ln_1_if_25_acc_nl[14:0];
  assign ln_1_if_25_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_25_acc_nl);
  assign nl_ln_1_if_24_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111000110101;
  assign ln_1_if_24_acc_nl = nl_ln_1_if_24_acc_nl[14:0];
  assign ln_1_if_24_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_24_acc_nl);
  assign nl_ln_1_if_23_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111100011001;
  assign ln_1_if_23_acc_nl = nl_ln_1_if_23_acc_nl[13:0];
  assign ln_1_if_23_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_23_acc_nl);
  assign nl_ln_1_if_22_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111000101111;
  assign ln_1_if_22_acc_nl = nl_ln_1_if_22_acc_nl[14:0];
  assign ln_1_if_22_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_22_acc_nl);
  assign nl_ln_1_if_21_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111110001011;
  assign ln_1_if_21_acc_nl = nl_ln_1_if_21_acc_nl[12:0];
  assign ln_1_if_21_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_21_acc_nl);
  assign nl_ln_1_if_20_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111000101001;
  assign ln_1_if_20_acc_nl = nl_ln_1_if_20_acc_nl[14:0];
  assign ln_1_if_20_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_20_acc_nl);
  assign nl_ln_1_if_19_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111100010011;
  assign ln_1_if_19_acc_nl = nl_ln_1_if_19_acc_nl[13:0];
  assign ln_1_if_19_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_19_acc_nl);
  assign nl_ln_1_if_18_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111000100011;
  assign ln_1_if_18_acc_nl = nl_ln_1_if_18_acc_nl[14:0];
  assign ln_1_if_18_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_18_acc_nl);
  assign nl_ln_1_if_17_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111000011111;
  assign ln_1_if_17_acc_nl = nl_ln_1_if_17_acc_nl[14:0];
  assign ln_1_if_17_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_17_acc_nl);
  assign nl_ln_1_if_16_acc_nl = conv_u2u_12_13(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:2])
      + 13'b1111110000111;
  assign ln_1_if_16_acc_nl = nl_ln_1_if_16_acc_nl[12:0];
  assign ln_1_if_16_acc_itm_12_1 = readslicef_13_1_12(ln_1_if_16_acc_nl);
  assign nl_ln_1_if_15_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111000011001;
  assign ln_1_if_15_acc_nl = nl_ln_1_if_15_acc_nl[14:0];
  assign ln_1_if_15_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_15_acc_nl);
  assign nl_ln_1_if_14_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111100001011;
  assign ln_1_if_14_acc_nl = nl_ln_1_if_14_acc_nl[13:0];
  assign ln_1_if_14_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_14_acc_nl);
  assign nl_ln_1_if_13_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111000010011;
  assign ln_1_if_13_acc_nl = nl_ln_1_if_13_acc_nl[14:0];
  assign ln_1_if_13_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_13_acc_nl);
  assign nl_ln_1_if_12_acc_nl = conv_u2u_10_11(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:4])
      + 11'b11111100001;
  assign ln_1_if_12_acc_nl = nl_ln_1_if_12_acc_nl[10:0];
  assign ln_1_if_12_acc_itm_10_1 = readslicef_11_1_10(ln_1_if_12_acc_nl);
  assign nl_ln_1_if_11_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111000001101;
  assign ln_1_if_11_acc_nl = nl_ln_1_if_11_acc_nl[14:0];
  assign ln_1_if_11_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_11_acc_nl);
  assign nl_ln_1_if_10_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111000001001;
  assign ln_1_if_10_acc_nl = nl_ln_1_if_10_acc_nl[14:0];
  assign ln_1_if_10_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_10_acc_nl);
  assign nl_ln_1_if_9_acc_nl = conv_u2u_13_14(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:1])
      + 14'b11111100000011;
  assign ln_1_if_9_acc_nl = nl_ln_1_if_9_acc_nl[13:0];
  assign ln_1_if_9_acc_itm_13_1 = readslicef_14_1_13(ln_1_if_9_acc_nl);
  assign nl_ln_1_if_8_acc_nl = conv_u2u_14_15(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1)
      + 15'b111111000000011;
  assign ln_1_if_8_acc_nl = nl_ln_1_if_8_acc_nl[14:0];
  assign ln_1_if_8_acc_itm_14_1 = readslicef_15_1_14(ln_1_if_8_acc_nl);
  assign nl_ln_1_if_4_acc_nl = conv_u2u_8_9(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:6])
      + 9'b111110101;
  assign ln_1_if_4_acc_nl = nl_ln_1_if_4_acc_nl[8:0];
  assign ln_1_if_4_acc_itm_8_1 = readslicef_9_1_8(ln_1_if_4_acc_nl);
  assign nl_ln_1_if_5_acc_nl = conv_u2u_7_8(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:7])
      + 8'b11111011;
  assign ln_1_if_5_acc_nl = nl_ln_1_if_5_acc_nl[7:0];
  assign ln_1_if_5_acc_itm_7_1 = readslicef_8_1_7(ln_1_if_5_acc_nl);
  assign nl_ln_1_if_3_acc_nl = conv_u2u_6_7(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:8])
      + 7'b1111101;
  assign ln_1_if_3_acc_nl = nl_ln_1_if_3_acc_nl[6:0];
  assign ln_1_if_3_acc_itm_6_1 = readslicef_7_1_6(ln_1_if_3_acc_nl);
  assign nl_ln_1_if_2_acc_nl = conv_u2u_8_9(operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1[13:6])
      + 9'b111110011;
  assign ln_1_if_2_acc_nl = nl_ln_1_if_2_acc_nl[8:0];
  assign ln_1_if_2_acc_itm_8_1 = readslicef_9_1_8(ln_1_if_2_acc_nl);
  assign if_4_for_1_and_stg_2_7_sva_1 = if_4_for_1_and_stg_1_3_sva_1 & (j_lpi_1_dfm_3_0_1[2]);
  assign if_4_for_1_and_stg_2_0_sva_1 = if_4_for_1_and_stg_1_0_sva_1 & (~ (j_lpi_1_dfm_3_0_1[2]));
  assign if_4_for_1_and_stg_2_6_sva_1 = if_4_for_1_and_stg_1_2_sva_1 & (j_lpi_1_dfm_3_0_1[2]);
  assign if_4_for_1_and_stg_2_1_sva_1 = if_4_for_1_and_stg_1_1_sva_1 & (~ (j_lpi_1_dfm_3_0_1[2]));
  assign if_4_for_1_and_stg_2_5_sva_1 = if_4_for_1_and_stg_1_1_sva_1 & (j_lpi_1_dfm_3_0_1[2]);
  assign if_4_for_1_and_stg_2_2_sva_1 = if_4_for_1_and_stg_1_2_sva_1 & (~ (j_lpi_1_dfm_3_0_1[2]));
  assign if_4_for_1_and_stg_2_4_sva_1 = if_4_for_1_and_stg_1_0_sva_1 & (j_lpi_1_dfm_3_0_1[2]);
  assign if_4_for_1_and_stg_2_3_sva_1 = if_4_for_1_and_stg_1_3_sva_1 & (~ (j_lpi_1_dfm_3_0_1[2]));
  assign if_4_for_1_and_stg_1_0_sva_1 = ~((j_lpi_1_dfm_3_0_1[1:0]!=2'b00));
  assign if_4_for_1_and_stg_1_1_sva_1 = (j_lpi_1_dfm_3_0_1[1:0]==2'b01);
  assign if_4_for_1_and_stg_1_2_sva_1 = (j_lpi_1_dfm_3_0_1[1:0]==2'b10);
  assign if_4_for_1_and_stg_1_3_sva_1 = (j_lpi_1_dfm_3_0_1[1:0]==2'b11);
  assign if_4_for_mux_50_tmp = MUX_v_10_2_2(asn_sft_lpi_1_dfm_st_1, count_sva, or_2_tmp);
  assign mux_3_tmp = MUX_v_2_2_2(reg_skip_ftd_1, skip_sva_1_1_0_1, or_324_cse);
  assign and_dcpl_24 = main_stage_0_2 & mux_1304_itm_1;
  assign and_dcpl_25 = (if_4_for_mux_50_tmp[9:8]==2'b11);
  assign and_dcpl_32 = (if_4_for_mux_50_tmp[1:0]==2'b11);
  assign nor_47_cse = ~(exitL_exit_if_4_for_2_lpi_1_dfm | exitL_exit_approx_sva);
  assign or_dcpl_1 = ~((~(((nor_47_cse & exit_if_4_for_lpi_1_dfm_2) | (j_1_3_0_sva_2[3]))
      & (if_4_for_1_acc_tmp[4]))) & nand_tmp);
  assign and_dcpl_39 = (if_4_for_mux_50_tmp[8:7]==2'b11);
  assign and_dcpl_41 = (if_4_for_mux_50_tmp[6:5]==2'b11);
  assign and_dcpl_42 = (if_4_for_mux_50_tmp[4:3]==2'b11);
  assign and_dcpl_43 = and_dcpl_42 & and_dcpl_41;
  assign or_dcpl_3 = or_2_tmp | (~ exit_if_4_for_lpi_1_dfm_2);
  assign and_dcpl_49 = (~(nand_112_cse & nand_tmp)) & and_dcpl_32 & or_dcpl_3 & (if_4_for_mux_50_tmp[2])
      & and_dcpl_43 & and_dcpl_39 & (if_4_for_mux_50_tmp[9]) & operator_24_14_false_AC_TRN_AC_WRAP_acc_itm_14_1;
  assign and_dcpl_59 = and_dcpl_32 & (if_4_for_mux_50_tmp[2]);
  assign and_dcpl_61 = or_dcpl_1 & and_dcpl_59 & and_dcpl_43 & and_dcpl_39 & (if_4_for_mux_50_tmp[9])
      & operator_24_14_false_AC_TRN_AC_WRAP_1_acc_itm_14_1;
  assign and_dcpl_66 = and_dcpl_59 & and_dcpl_42 & and_dcpl_41 & (if_4_for_mux_50_tmp[7])
      & and_dcpl_25;
  assign and_dcpl_67 = ~((((~(exitL_exit_if_4_for_2_lpi_1_dfm | (~ exit_if_4_for_lpi_1_dfm_2)
      | exitL_exit_approx_sva)) | (j_1_3_0_sva_2[3])) & (if_4_for_1_acc_tmp[4]))
      | nand_tmp);
  assign or_dcpl_10 = ~(main_stage_0_3 & mux_1304_itm_2);
  assign or_dcpl_14 = ~((asn_sft_lpi_1_dfm_st_1[4:2]==3'b111));
  assign or_dcpl_20 = (~((asn_sft_lpi_1_dfm_st_1[0]) & (asn_sft_lpi_1_dfm_st_1[9])
      & (asn_sft_lpi_1_dfm_st_1[8]))) | (~((asn_sft_lpi_1_dfm_st_1[7:5]==3'b111)));
  assign or_dcpl_26 = shift_reg_1_sva_1 | shift_reg_1_sva_0;
  assign or_dcpl_27 = (mux_3_tmp[0]) | shift_reg_1_sva_2;
  assign or_dcpl_28 = or_dcpl_27 | or_dcpl_26;
  assign or_dcpl_29 = epsilon_rsci_idat | (mux_3_tmp[1]);
  assign mux_tmp_4 = MUX_s_1_2_2((~ exitL_exit_if_4_for_2_lpi_1_dfm), epsilon_rsci_idat,
      exitL_exit_approx_sva);
  assign or_dcpl_33 = (mux_3_tmp[0]) | (~ shift_reg_1_sva_2);
  assign or_dcpl_34 = or_dcpl_33 | or_dcpl_26;
  assign or_dcpl_37 = (~ epsilon_rsci_idat) | (mux_3_tmp[1]);
  assign mux_1310_itm = MUX_s_1_2_2(exitL_exit_if_4_for_2_lpi_1_dfm, epsilon_rsci_idat,
      exitL_exit_approx_sva);
  assign or_dcpl_43 = shift_reg_1_sva_1 | (~ shift_reg_1_sva_0);
  assign or_dcpl_44 = or_dcpl_27 | or_dcpl_43;
  assign or_dcpl_47 = or_dcpl_33 | or_dcpl_43;
  assign or_dcpl_54 = (~ shift_reg_1_sva_1) | shift_reg_1_sva_0;
  assign or_dcpl_55 = or_dcpl_33 | or_dcpl_54;
  assign or_dcpl_58 = or_dcpl_27 | or_dcpl_54;
  assign or_dcpl_65 = ~(shift_reg_1_sva_1 & shift_reg_1_sva_0);
  assign or_dcpl_66 = or_dcpl_33 | or_dcpl_65;
  assign or_dcpl_69 = or_dcpl_27 | or_dcpl_65;
  assign or_dcpl_76 = (mux_3_tmp[1]) | shift_reg_1_sva_1;
  assign or_dcpl_77 = or_dcpl_76 | shift_reg_1_sva_0;
  assign or_dcpl_80 = (mux_3_tmp[1]) | (~ shift_reg_1_sva_1);
  assign or_dcpl_81 = or_dcpl_80 | shift_reg_1_sva_0;
  assign or_dcpl_88 = or_dcpl_76 | (~ shift_reg_1_sva_0);
  assign or_dcpl_91 = or_dcpl_80 | (~ shift_reg_1_sva_0);
  assign or_dcpl_98 = epsilon_rsci_idat | (~ shift_reg_1_sva_0);
  assign or_tmp_12 = shift_reg_1_sva_1 | shift_reg_1_sva_2 | (~ first_sva) | (mux_3_tmp!=2'b00);
  assign or_tmp_14 = saved_reg_sva_2 | (~ or_247_cse);
  assign mux_tmp_9 = MUX_s_1_2_2((~ or_226_cse), or_222_cse, saved_reg_sva_2);
  assign mux_1315_nl = MUX_s_1_2_2(mux_tmp_9, or_tmp_14, shift_reg_1_sva_1);
  assign mux_tmp_11 = MUX_s_1_2_2(mux_1315_nl, or_tmp_12, saved_reg_sva_1);
  assign or_dcpl_100 = saved_reg_sva_2 | saved_reg_sva_1;
  assign or_dcpl_102 = (~ or_247_cse) | epsilon_rsci_idat;
  assign or_dcpl_104 = epsilon_rsci_idat | shift_reg_1_sva_0;
  assign or_tmp_19 = (~ shift_reg_1_sva_1) | shift_reg_1_sva_2 | (~ first_sva) |
      (mux_3_tmp!=2'b00);
  assign mux_1320_nl = MUX_s_1_2_2(or_tmp_14, mux_tmp_9, shift_reg_1_sva_1);
  assign mux_tmp_16 = MUX_s_1_2_2(or_tmp_19, mux_1320_nl, saved_reg_sva_1);
  assign or_tmp_21 = (~ saved_reg_sva_2) | saved_reg_sva_1;
  assign and_tmp = shift_reg_1_sva_1 & epsilon_rsci_idat;
  assign or_tmp_27 = shift_reg_1_sva_1 | (~ shift_reg_1_sva_2) | (~ first_sva) |
      (mux_3_tmp!=2'b00);
  assign and_tmp_1 = saved_reg_sva_2 & or_247_cse;
  assign mux_1326_nl = MUX_s_1_2_2(mux_tmp_9, and_tmp_1, shift_reg_1_sva_1);
  assign mux_tmp_22 = MUX_s_1_2_2((~ mux_1326_nl), or_tmp_27, saved_reg_sva_1);
  assign mux_tmp_23 = MUX_s_1_2_2(or_226_cse, or_222_cse, shift_reg_1_sva_1);
  assign mux_tmp_24 = MUX_s_1_2_2((~ or_222_cse), or_226_cse, saved_reg_sva_2);
  assign nor_tmp_5 = saved_reg_sva_2 & saved_reg_sva_1;
  assign or_tmp_29 = (~ shift_reg_1_sva_1) | (~ shift_reg_1_sva_2) | (~ first_sva)
      | (mux_3_tmp!=2'b00);
  assign mux_1335_nl = MUX_s_1_2_2(and_tmp_1, mux_tmp_9, shift_reg_1_sva_1);
  assign not_tmp_48 = MUX_s_1_2_2(or_tmp_29, (~ mux_1335_nl), saved_reg_sva_1);
  assign or_dcpl_118 = ~(epsilon_rsci_idat & shift_reg_1_sva_0);
  assign or_dcpl_121 = (~ epsilon_rsci_idat) | shift_reg_1_sva_0;
  assign or_dcpl_132 = ~(or_247_cse & epsilon_rsci_idat);
  assign or_dcpl_139 = (~ epsilon_rsci_idat) | or_dcpl_65;
  assign or_dcpl_144 = epsilon_rsci_idat | or_dcpl_26;
  assign mux_1356_nl = MUX_s_1_2_2((~ or_247_cse), or_247_cse, epsilon_rsci_idat);
  assign mux_tmp_53 = MUX_s_1_2_2((~ or_247_cse), mux_1356_nl, exitL_exit_approx_sva);
  assign or_209_nl = (~ epsilon_rsci_idat) | (~ first_sva) | (mux_3_tmp!=2'b00);
  assign mux_1361_nl = MUX_s_1_2_2(or_247_cse, or_209_nl, exitL_exit_approx_sva);
  assign or_207_nl = epsilon_rsci_idat | (~ first_sva) | (mux_3_tmp!=2'b00);
  assign mux_1360_nl = MUX_s_1_2_2(or_247_cse, or_207_nl, exitL_exit_approx_sva);
  assign mux_tmp_57 = MUX_s_1_2_2(mux_1361_nl, mux_1360_nl, shift_reg_1_sva_2);
  assign or_dcpl_151 = epsilon_rsci_idat | or_dcpl_65;
  assign or_dcpl_154 = (~ epsilon_rsci_idat) | or_dcpl_26;
  assign mux_tmp_61 = MUX_s_1_2_2(nor_63_cse, or_222_cse, saved_reg_sva_2);
  assign or_dcpl_164 = epsilon_rsci_idat | or_dcpl_43;
  assign or_dcpl_170 = epsilon_rsci_idat | or_dcpl_54;
  assign or_dcpl_174 = (~ epsilon_rsci_idat) | or_dcpl_43;
  assign or_dcpl_180 = or_247_cse | nor_47_cse;
  assign or_dcpl_185 = ~((if_4_for_mux_50_tmp[4:3]==2'b11));
  assign or_dcpl_188 = ~((if_4_for_mux_50_tmp[2:0]==3'b111));
  assign or_tmp_82 = saved_reg_sva_0 | saved_reg_sva_1 | saved_reg_sva_2;
  assign or_tmp_83 = or_tmp_82 | (~ and_276_cse);
  assign or_tmp_85 = or_dcpl_100 | (~ and_276_cse);
  assign not_tmp_87 = ~(shift_reg_1_sva_1 & (count_sva==10'b1111111111));
  assign or_tmp_86 = saved_reg_sva_2 | not_tmp_87;
  assign mux_1408_nl = MUX_s_1_2_2(or_tmp_86, or_tmp_85, shift_reg_1_sva_0);
  assign mux_tmp_96 = MUX_s_1_2_2(mux_1408_nl, or_tmp_83, epsilon_rsci_idat);
  assign or_tmp_88 = first_sva | saved_reg_sva_0 | saved_reg_sva_1 | saved_reg_sva_2
      | (~ and_276_cse);
  assign or_tmp_89 = shift_reg_1_sva_2 | shift_reg_1_sva_1;
  assign or_tmp_90 = or_tmp_89 | (~ and_276_cse);
  assign not_tmp_88 = shift_reg_1_sva_1 & (~ and_276_cse);
  assign mux_1414_nl = MUX_s_1_2_2(not_tmp_88, shift_reg_1_sva_1, saved_reg_sva_2);
  assign mux_1415_nl = MUX_s_1_2_2(or_tmp_86, mux_1414_nl, shift_reg_1_sva_2);
  assign mux_1413_nl = MUX_s_1_2_2(not_tmp_87, shift_reg_1_sva_1, shift_reg_1_sva_2);
  assign mux_1416_nl = MUX_s_1_2_2(mux_1415_nl, mux_1413_nl, first_sva);
  assign mux_1412_nl = MUX_s_1_2_2(or_tmp_85, or_tmp_90, first_sva);
  assign mux_tmp_104 = MUX_s_1_2_2(mux_1416_nl, mux_1412_nl, shift_reg_1_sva_0);
  assign mux_1410_nl = MUX_s_1_2_2(or_tmp_83, or_tmp_90, first_sva);
  assign mux_1411_nl = MUX_s_1_2_2(mux_1410_nl, or_tmp_88, shift_reg_1_sva_0);
  assign mux_tmp_105 = MUX_s_1_2_2(mux_tmp_104, mux_1411_nl, epsilon_rsci_idat);
  assign or_tmp_93 = shift_reg_1_sva_1 | and_276_cse;
  assign or_327_cse = shift_reg_1_sva_1 | (~ and_276_cse);
  assign mux_1422_nl = MUX_s_1_2_2(not_tmp_88, or_tmp_93, or_tmp_82);
  assign mux_1423_nl = MUX_s_1_2_2(or_tmp_83, mux_1422_nl, shift_reg_1_sva_2);
  assign mux_1421_nl = MUX_s_1_2_2(or_327_cse, or_tmp_93, shift_reg_1_sva_2);
  assign mux_1424_nl = MUX_s_1_2_2(mux_1423_nl, mux_1421_nl, first_sva);
  assign mux_1425_nl = MUX_s_1_2_2(mux_1424_nl, or_tmp_88, shift_reg_1_sva_0);
  assign mux_tmp_113 = MUX_s_1_2_2(mux_tmp_104, mux_1425_nl, epsilon_rsci_idat);
  assign not_tmp_91 = ~((count_sva==10'b1111111111));
  assign or_tmp_100 = epsilon_rsci_idat | not_tmp_91;
  assign not_tmp_92 = ~(saved_reg_sva_0 & epsilon_rsci_idat & (count_sva==10'b1111111111));
  assign mux_1431_nl = MUX_s_1_2_2(not_tmp_92, or_tmp_100, saved_reg_sva_1);
  assign or_tmp_101 = saved_reg_sva_2 | mux_1431_nl;
  assign or_335_nl = saved_reg_sva_1 | not_tmp_92;
  assign mux_tmp_119 = MUX_s_1_2_2(or_335_nl, or_tmp_100, saved_reg_sva_2);
  assign or_tmp_104 = or_dcpl_100 | not_tmp_92;
  assign mux_1434_nl = MUX_s_1_2_2(or_tmp_104, or_tmp_101, shift_reg_1_sva_0);
  assign mux_1433_nl = MUX_s_1_2_2(mux_tmp_119, or_tmp_101, shift_reg_1_sva_0);
  assign mux_tmp_122 = MUX_s_1_2_2(mux_1434_nl, mux_1433_nl, shift_reg_1_sva_1);
  assign or_tmp_105 = shift_reg_1_sva_2 | epsilon_rsci_idat;
  assign or_341_cse = (~ shift_reg_1_sva_2) | epsilon_rsci_idat | not_tmp_91;
  assign mux_1437_nl = MUX_s_1_2_2(mux_tmp_119, or_341_cse, first_sva);
  assign or_339_nl = or_tmp_105 | not_tmp_91;
  assign mux_1436_nl = MUX_s_1_2_2(or_tmp_101, or_339_nl, first_sva);
  assign mux_tmp_125 = MUX_s_1_2_2(mux_1437_nl, mux_1436_nl, shift_reg_1_sva_0);
  assign nand_116_cse = ~(epsilon_rsci_idat & (count_sva==10'b1111111111));
  assign or_342_nl = shift_reg_1_sva_2 | nand_116_cse;
  assign mux_tmp_126 = MUX_s_1_2_2(or_tmp_101, or_342_nl, first_sva);
  assign mux_1440_nl = MUX_s_1_2_2(or_tmp_104, (~ epsilon_rsci_idat), shift_reg_1_sva_2);
  assign nand_117_nl = ~(shift_reg_1_sva_2 & epsilon_rsci_idat);
  assign mux_1441_nl = MUX_s_1_2_2(mux_1440_nl, nand_117_nl, first_sva);
  assign mux_1442_nl = MUX_s_1_2_2(mux_1441_nl, mux_tmp_126, shift_reg_1_sva_0);
  assign mux_tmp_130 = MUX_s_1_2_2(mux_1442_nl, mux_tmp_125, shift_reg_1_sva_1);
  assign mux_1446_nl = MUX_s_1_2_2(or_tmp_104, (~ or_tmp_100), shift_reg_1_sva_2);
  assign nand_118_nl = ~(shift_reg_1_sva_2 & or_tmp_100);
  assign mux_1447_nl = MUX_s_1_2_2(mux_1446_nl, nand_118_nl, first_sva);
  assign mux_1448_nl = MUX_s_1_2_2(mux_1447_nl, mux_tmp_126, shift_reg_1_sva_0);
  assign mux_tmp_136 = MUX_s_1_2_2(mux_1448_nl, mux_tmp_125, shift_reg_1_sva_1);
  assign or_350_nl = shift_reg_1_sva_2 | shift_reg_1_sva_1 | shift_reg_1_sva_0;
  assign or_349_nl = (skip_sva_1_1_0_1!=2'b00) | shift_reg_1_sva_2 | shift_reg_1_sva_1
      | shift_reg_1_sva_0;
  assign mux_tmp_141 = MUX_s_1_2_2(or_350_nl, or_349_nl, or_324_cse);
  assign mux_1455_nl = MUX_s_1_2_2((~ saved_reg_sva_0), shift_reg_1_sva_0, saved_reg_sva_1);
  assign mux_tmp_143 = MUX_s_1_2_2(mux_1455_nl, or_dcpl_26, saved_reg_sva_2);
  assign mux_1457_nl = MUX_s_1_2_2((~ shift_reg_1_sva_0), shift_reg_1_sva_0, shift_reg_1_sva_1);
  assign mux_tmp_145 = MUX_s_1_2_2(mux_1457_nl, or_dcpl_26, shift_reg_1_sva_2);
  assign or_tmp_121 = ~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_lpi_1_dfm_1_3_0==4'b0001));
  assign or_tmp_125 = saved_reg_sva_0 | (~ saved_reg_sva_1) | saved_reg_sva_2 | (~
      and_276_cse);
  assign not_tmp_104 = ~(saved_reg_sva_2 & (count_sva==10'b1111111111));
  assign or_tmp_127 = saved_reg_sva_2 | (~ and_276_cse);
  assign mux_1468_nl = MUX_s_1_2_2(or_tmp_125, or_tmp_127, shift_reg_1_sva_1);
  assign nand_71_nl = ~(epsilon_rsci_idat & (~ mux_1468_nl));
  assign or_359_nl = saved_reg_sva_1 | not_tmp_104;
  assign mux_1467_nl = MUX_s_1_2_2(or_359_nl, or_tmp_125, epsilon_rsci_idat);
  assign mux_tmp_156 = MUX_s_1_2_2(nand_71_nl, mux_1467_nl, shift_reg_1_sva_0);
  assign or_tmp_129 = first_sva | saved_reg_sva_0 | (~ saved_reg_sva_1) | saved_reg_sva_2
      | (~ and_276_cse);
  assign or_tmp_131 = first_sva | saved_reg_sva_1 | not_tmp_104;
  assign nor_189_nl = ~(shift_reg_1_sva_2 | (~ or_tmp_131));
  assign mux_tmp_157 = MUX_s_1_2_2(nor_189_nl, or_tmp_131, shift_reg_1_sva_1);
  assign or_tmp_133 = first_sva | saved_reg_sva_2;
  assign mux_1472_nl = MUX_s_1_2_2(or_tmp_127, (~ and_276_cse), first_sva);
  assign or_367_nl = or_tmp_133 | (~ and_276_cse);
  assign mux_1473_nl = MUX_s_1_2_2(mux_1472_nl, or_367_nl, shift_reg_1_sva_2);
  assign mux_1474_nl = MUX_s_1_2_2(or_tmp_129, mux_1473_nl, shift_reg_1_sva_1);
  assign nand_tmp_13 = ~(epsilon_rsci_idat & (~ mux_1474_nl));
  assign mux_1471_nl = MUX_s_1_2_2(mux_tmp_157, or_tmp_129, epsilon_rsci_idat);
  assign mux_tmp_162 = MUX_s_1_2_2(nand_tmp_13, mux_1471_nl, shift_reg_1_sva_0);
  assign nor_87_cse = ~(shift_reg_1_sva_1 | (~ shift_reg_1_sva_2));
  assign and_308_nl = (first_sva | saved_reg_sva_0 | (~ saved_reg_sva_1) | saved_reg_sva_2)
      & (count_sva==10'b1111111111);
  assign mux_1478_nl = MUX_s_1_2_2(or_tmp_129, and_308_nl, nor_87_cse);
  assign mux_1479_nl = MUX_s_1_2_2(mux_tmp_157, mux_1478_nl, epsilon_rsci_idat);
  assign mux_tmp_167 = MUX_s_1_2_2(nand_tmp_13, mux_1479_nl, shift_reg_1_sva_0);
  assign or_tmp_143 = epsilon_rsci_idat | (~ saved_reg_sva_1) | saved_reg_sva_0 |
      saved_reg_sva_2 | not_tmp_91;
  assign or_378_nl = saved_reg_sva_0 | saved_reg_sva_2 | not_tmp_91;
  assign mux_tmp_172 = MUX_s_1_2_2(not_tmp_104, or_378_nl, saved_reg_sva_1);
  assign or_tmp_146 = epsilon_rsci_idat | mux_tmp_172;
  assign mux_tmp_173 = MUX_s_1_2_2(or_tmp_146, or_tmp_143, shift_reg_1_sva_0);
  assign or_380_nl = saved_reg_sva_2 | not_tmp_91;
  assign mux_tmp_174 = MUX_s_1_2_2(mux_tmp_172, or_380_nl, epsilon_rsci_idat);
  assign or_382_nl = shift_reg_1_sva_0 | shift_reg_1_sva_2 | epsilon_rsci_idat |
      not_tmp_91;
  assign mux_tmp_177 = MUX_s_1_2_2(mux_tmp_173, or_382_nl, first_sva);
  assign mux_1493_nl = MUX_s_1_2_2(epsilon_rsci_idat, or_tmp_143, shift_reg_1_sva_2);
  assign mux_1494_nl = MUX_s_1_2_2(mux_tmp_174, mux_1493_nl, shift_reg_1_sva_0);
  assign mux_1491_nl = MUX_s_1_2_2((~ and_294_cse), or_tmp_100, shift_reg_1_sva_2);
  assign mux_1492_nl = MUX_s_1_2_2(mux_1491_nl, or_tmp_105, shift_reg_1_sva_0);
  assign mux_1495_nl = MUX_s_1_2_2(mux_1494_nl, mux_1492_nl, first_sva);
  assign mux_tmp_183 = MUX_s_1_2_2(mux_1495_nl, mux_tmp_177, shift_reg_1_sva_1);
  assign mux_tmp_186 = MUX_s_1_2_2(mux_tmp_174, or_tmp_146, shift_reg_1_sva_2);
  assign or_387_cse = shift_reg_1_sva_2 | and_294_cse;
  assign mux_1503_nl = MUX_s_1_2_2(and_294_cse, or_tmp_143, shift_reg_1_sva_2);
  assign mux_1504_nl = MUX_s_1_2_2(mux_tmp_186, mux_1503_nl, shift_reg_1_sva_0);
  assign nand_123_nl = ~((shift_reg_1_sva_2 | epsilon_rsci_idat | saved_reg_sva_2)
      & (count_sva==10'b1111111111));
  assign mux_1502_nl = MUX_s_1_2_2(nand_123_nl, or_387_cse, shift_reg_1_sva_0);
  assign mux_1505_nl = MUX_s_1_2_2(mux_1504_nl, mux_1502_nl, first_sva);
  assign mux_tmp_193 = MUX_s_1_2_2(mux_1505_nl, mux_tmp_177, shift_reg_1_sva_1);
  assign nor_tmp_32 = saved_reg_sva_1 & saved_reg_sva_0 & (count_sva==10'b1111111111);
  assign or_393_nl = (~ shift_reg_1_sva_1) | shift_reg_1_sva_0 | (~ and_276_cse);
  assign mux_tmp_198 = MUX_s_1_2_2((~ nor_tmp_32), or_393_nl, saved_reg_sva_2);
  assign not_tmp_120 = ~(saved_reg_sva_2 & saved_reg_sva_1 & shift_reg_1_sva_0 &
      (count_sva==10'b1111111111));
  assign mux_tmp_199 = MUX_s_1_2_2(not_tmp_120, mux_tmp_198, epsilon_rsci_idat);
  assign or_tmp_161 = shift_reg_1_sva_0 | (~ and_276_cse);
  assign mux_tmp_200 = MUX_s_1_2_2((~ shift_reg_1_sva_0), or_tmp_161, shift_reg_1_sva_1);
  assign nor_tmp_35 = epsilon_rsci_idat & shift_reg_1_sva_1 & shift_reg_1_sva_0 &
      (count_sva==10'b1111111111);
  assign and_317_cse = saved_reg_sva_0 & (count_sva==10'b1111111111);
  assign or_395_nl = shift_reg_1_sva_0 | and_317_cse;
  assign mux_1516_nl = MUX_s_1_2_2(shift_reg_1_sva_0, or_395_nl, saved_reg_sva_1);
  assign mux_1517_nl = MUX_s_1_2_2(mux_1516_nl, nor_tmp_32, shift_reg_1_sva_1);
  assign mux_tmp_205 = MUX_s_1_2_2((~ mux_1517_nl), mux_tmp_200, saved_reg_sva_2);
  assign nand_125_cse = ~(shift_reg_1_sva_1 & shift_reg_1_sva_0 & (count_sva==10'b1111111111));
  assign mux_1519_nl = MUX_s_1_2_2(not_tmp_120, mux_tmp_205, epsilon_rsci_idat);
  assign mux_1520_nl = MUX_s_1_2_2(mux_tmp_199, mux_1519_nl, shift_reg_1_sva_2);
  assign mux_1514_nl = MUX_s_1_2_2(nand_125_cse, mux_tmp_200, epsilon_rsci_idat);
  assign mux_1515_nl = MUX_s_1_2_2((~ nor_tmp_35), mux_1514_nl, shift_reg_1_sva_2);
  assign mux_tmp_208 = MUX_s_1_2_2(mux_1520_nl, mux_1515_nl, first_sva);
  assign mux_tmp_211 = MUX_s_1_2_2((~ or_tmp_161), and_276_cse, saved_reg_sva_1);
  assign and_319_nl = saved_reg_sva_1 & shift_reg_1_sva_0 & (count_sva==10'b1111111111);
  assign mux_1525_nl = MUX_s_1_2_2(and_319_nl, mux_tmp_211, shift_reg_1_sva_1);
  assign nand_126_nl = ~(saved_reg_sva_2 & mux_1525_nl);
  assign mux_tmp_213 = MUX_s_1_2_2(nand_126_nl, mux_tmp_198, epsilon_rsci_idat);
  assign not_tmp_127 = shift_reg_1_sva_0 & (~ and_276_cse);
  assign nor_192_nl = ~(shift_reg_1_sva_1 | (~ shift_reg_1_sva_0) | and_276_cse);
  assign mux_1531_nl = MUX_s_1_2_2(not_tmp_127, shift_reg_1_sva_0, saved_reg_sva_1);
  assign mux_1532_nl = MUX_s_1_2_2(mux_1531_nl, mux_tmp_211, shift_reg_1_sva_1);
  assign mux_1533_nl = MUX_s_1_2_2(nor_192_nl, mux_1532_nl, saved_reg_sva_2);
  assign mux_1534_nl = MUX_s_1_2_2((~ mux_1533_nl), mux_tmp_205, epsilon_rsci_idat);
  assign mux_1535_nl = MUX_s_1_2_2(mux_tmp_213, mux_1534_nl, shift_reg_1_sva_2);
  assign mux_1528_nl = MUX_s_1_2_2(not_tmp_127, and_276_cse, shift_reg_1_sva_1);
  assign mux_1527_nl = MUX_s_1_2_2(shift_reg_1_sva_0, and_276_cse, shift_reg_1_sva_1);
  assign mux_1529_nl = MUX_s_1_2_2(mux_1528_nl, mux_1527_nl, epsilon_rsci_idat);
  assign mux_1530_nl = MUX_s_1_2_2(nor_tmp_35, mux_1529_nl, shift_reg_1_sva_2);
  assign not_tmp_131 = MUX_s_1_2_2(mux_1535_nl, (~ mux_1530_nl), first_sva);
  assign or_tmp_170 = shift_reg_1_sva_1 | (~ saved_reg_sva_2) | shift_reg_1_sva_0
      | (~ and_276_cse);
  assign not_tmp_135 = ~(saved_reg_sva_0 & saved_reg_sva_1 & (count_sva==10'b1111111111));
  assign or_405_nl = (~ saved_reg_sva_1) | shift_reg_1_sva_0 | (~ and_276_cse);
  assign mux_tmp_228 = MUX_s_1_2_2(not_tmp_135, or_405_nl, saved_reg_sva_2);
  assign or_tmp_176 = shift_reg_1_sva_0 | and_276_cse;
  assign mux_1544_nl = MUX_s_1_2_2(shift_reg_1_sva_0, or_tmp_176, saved_reg_sva_2);
  assign or_408_nl = (~ saved_reg_sva_2) | shift_reg_1_sva_0 | (~ and_276_cse);
  assign mux_1545_nl = MUX_s_1_2_2((~ mux_1544_nl), or_408_nl, shift_reg_1_sva_2);
  assign mux_1543_nl = MUX_s_1_2_2((~ shift_reg_1_sva_0), or_tmp_161, shift_reg_1_sva_2);
  assign mux_tmp_233 = MUX_s_1_2_2(mux_1545_nl, mux_1543_nl, first_sva);
  assign nand_128_cse = ~(shift_reg_1_sva_0 & (count_sva==10'b1111111111));
  assign mux_1547_cse = MUX_s_1_2_2(nand_128_cse, or_tmp_161, shift_reg_1_sva_2);
  assign mux_tmp_235 = MUX_s_1_2_2(mux_tmp_228, mux_1547_cse, first_sva);
  assign or_411_nl = first_sva | mux_tmp_228;
  assign mux_1549_nl = MUX_s_1_2_2(or_411_nl, mux_tmp_235, shift_reg_1_sva_1);
  assign or_410_nl = shift_reg_1_sva_1 | mux_tmp_233;
  assign mux_tmp_237 = MUX_s_1_2_2(mux_1549_nl, or_410_nl, epsilon_rsci_idat);
  assign mux_tmp_240 = MUX_s_1_2_2(not_tmp_135, or_tmp_161, saved_reg_sva_2);
  assign nand_tmp_16 = ~(shift_reg_1_sva_0 & (~ and_276_cse));
  assign mux_1558_cse = MUX_s_1_2_2((~ and_276_cse), and_276_cse, shift_reg_1_sva_0);
  assign and_324_nl = saved_reg_sva_0 & saved_reg_sva_1;
  assign mux_1559_nl = MUX_s_1_2_2(nand_tmp_16, (~ or_tmp_176), and_324_nl);
  assign mux_1560_nl = MUX_s_1_2_2(mux_1559_nl, mux_1558_cse, saved_reg_sva_2);
  assign mux_1561_nl = MUX_s_1_2_2(mux_1560_nl, mux_tmp_240, shift_reg_1_sva_2);
  assign mux_1557_nl = MUX_s_1_2_2(nand_tmp_16, or_tmp_161, shift_reg_1_sva_2);
  assign mux_1562_nl = MUX_s_1_2_2(mux_1561_nl, mux_1557_nl, first_sva);
  assign mux_1563_nl = MUX_s_1_2_2(mux_1562_nl, mux_tmp_235, shift_reg_1_sva_1);
  assign nand_129_nl = ~(first_sva & shift_reg_1_sva_2 & (~ shift_reg_1_sva_0) &
      and_276_cse);
  assign mux_1556_nl = MUX_s_1_2_2(mux_tmp_233, nand_129_nl, shift_reg_1_sva_1);
  assign mux_tmp_251 = MUX_s_1_2_2(mux_1563_nl, mux_1556_nl, epsilon_rsci_idat);
  assign or_tmp_186 = saved_reg_sva_0 | saved_reg_sva_1;
  assign or_tmp_187 = or_tmp_186 | (~ and_276_cse);
  assign or_421_nl = saved_reg_sva_1 | nand_128_cse;
  assign mux_tmp_256 = MUX_s_1_2_2(or_421_nl, or_tmp_187, saved_reg_sva_2);
  assign or_tmp_190 = (~ shift_reg_1_sva_1) | saved_reg_sva_2 | nand_128_cse;
  assign mux_tmp_259 = MUX_s_1_2_2(mux_tmp_256, mux_1547_cse, first_sva);
  assign or_426_nl = saved_reg_sva_2 | nand_128_cse;
  assign mux_1575_nl = MUX_s_1_2_2(not_tmp_127, shift_reg_1_sva_0, saved_reg_sva_2);
  assign mux_1576_nl = MUX_s_1_2_2(or_426_nl, mux_1575_nl, shift_reg_1_sva_2);
  assign mux_1574_nl = MUX_s_1_2_2(nand_128_cse, shift_reg_1_sva_0, shift_reg_1_sva_2);
  assign mux_tmp_264 = MUX_s_1_2_2(mux_1576_nl, mux_1574_nl, first_sva);
  assign nand_77_nl = ~(shift_reg_1_sva_1 & (~ mux_tmp_264));
  assign or_424_nl = first_sva | mux_tmp_256;
  assign mux_1573_nl = MUX_s_1_2_2(mux_tmp_259, or_424_nl, shift_reg_1_sva_1);
  assign mux_tmp_265 = MUX_s_1_2_2(nand_77_nl, mux_1573_nl, epsilon_rsci_idat);
  assign mux_tmp_268 = MUX_s_1_2_2(nand_128_cse, or_tmp_187, saved_reg_sva_2);
  assign or_432_nl = (~ first_sva) | shift_reg_1_sva_2 | nand_128_cse;
  assign mux_1591_nl = MUX_s_1_2_2(or_432_nl, mux_tmp_264, shift_reg_1_sva_1);
  assign mux_1586_nl = MUX_s_1_2_2(and_276_cse, (~ and_276_cse), shift_reg_1_sva_0);
  assign mux_1585_nl = MUX_s_1_2_2(not_tmp_127, or_tmp_176, or_tmp_186);
  assign mux_1587_nl = MUX_s_1_2_2(mux_1586_nl, mux_1585_nl, saved_reg_sva_2);
  assign mux_1588_nl = MUX_s_1_2_2(mux_tmp_268, mux_1587_nl, shift_reg_1_sva_2);
  assign mux_1584_nl = MUX_s_1_2_2(nand_128_cse, or_tmp_176, shift_reg_1_sva_2);
  assign mux_1589_nl = MUX_s_1_2_2(mux_1588_nl, mux_1584_nl, first_sva);
  assign mux_1590_nl = MUX_s_1_2_2(mux_tmp_259, mux_1589_nl, shift_reg_1_sva_1);
  assign mux_tmp_279 = MUX_s_1_2_2(mux_1591_nl, mux_1590_nl, epsilon_rsci_idat);
  assign or_tmp_205 = saved_reg_sva_2 | saved_reg_sva_1 | shift_reg_1_sva_0 | (~
      and_276_cse);
  assign or_441_nl = shift_reg_1_sva_1 | nand_128_cse;
  assign mux_tmp_284 = MUX_s_1_2_2(or_441_nl, or_tmp_187, saved_reg_sva_2);
  assign mux_tmp_285 = MUX_s_1_2_2(mux_tmp_284, or_tmp_205, epsilon_rsci_idat);
  assign or_tmp_209 = epsilon_rsci_idat | shift_reg_1_sva_1 | shift_reg_1_sva_0;
  assign or_tmp_210 = or_tmp_209 | (~ and_276_cse);
  assign mux_tmp_286 = MUX_s_1_2_2(nand_128_cse, shift_reg_1_sva_0, shift_reg_1_sva_1);
  assign or_446_cse = saved_reg_sva_0 | (~ and_276_cse);
  assign and_255_nl = shift_reg_1_sva_0 & or_446_cse;
  assign mux_1602_nl = MUX_s_1_2_2(and_255_nl, shift_reg_1_sva_0, saved_reg_sva_1);
  assign mux_1603_nl = MUX_s_1_2_2(or_tmp_187, mux_1602_nl, shift_reg_1_sva_1);
  assign mux_tmp_291 = MUX_s_1_2_2(mux_tmp_286, mux_1603_nl, saved_reg_sva_2);
  assign mux_1605_nl = MUX_s_1_2_2(mux_tmp_291, or_tmp_205, epsilon_rsci_idat);
  assign mux_1606_nl = MUX_s_1_2_2(mux_1605_nl, mux_tmp_285, shift_reg_1_sva_2);
  assign or_445_nl = or_dcpl_26 | (~ and_276_cse);
  assign mux_1600_nl = MUX_s_1_2_2(mux_tmp_286, or_445_nl, epsilon_rsci_idat);
  assign mux_1601_nl = MUX_s_1_2_2(mux_1600_nl, or_tmp_210, shift_reg_1_sva_2);
  assign mux_tmp_294 = MUX_s_1_2_2(mux_1606_nl, mux_1601_nl, first_sva);
  assign or_tmp_216 = saved_reg_sva_1 | shift_reg_1_sva_0;
  assign not_tmp_151 = ~(((~ saved_reg_sva_1) | shift_reg_1_sva_0) & (count_sva==10'b1111111111));
  assign or_450_nl = or_tmp_216 | (~ and_276_cse);
  assign mux_1610_nl = MUX_s_1_2_2(not_tmp_151, or_450_nl, shift_reg_1_sva_1);
  assign or_452_nl = saved_reg_sva_2 | mux_1610_nl;
  assign mux_tmp_298 = MUX_s_1_2_2(mux_tmp_284, or_452_nl, epsilon_rsci_idat);
  assign mux_1616_nl = MUX_s_1_2_2(shift_reg_1_sva_0, or_tmp_176, saved_reg_sva_1);
  assign mux_1617_nl = MUX_s_1_2_2(not_tmp_151, mux_1616_nl, shift_reg_1_sva_1);
  assign or_455_nl = (~ shift_reg_1_sva_1) | shift_reg_1_sva_0 | and_276_cse;
  assign mux_1618_nl = MUX_s_1_2_2(mux_1617_nl, or_455_nl, saved_reg_sva_2);
  assign mux_1619_nl = MUX_s_1_2_2(mux_tmp_291, mux_1618_nl, epsilon_rsci_idat);
  assign mux_1620_nl = MUX_s_1_2_2(mux_1619_nl, mux_tmp_298, shift_reg_1_sva_2);
  assign mux_1613_nl = MUX_s_1_2_2((~ and_276_cse), shift_reg_1_sva_0, shift_reg_1_sva_1);
  assign mux_1612_nl = MUX_s_1_2_2((~ and_276_cse), or_tmp_176, shift_reg_1_sva_1);
  assign mux_1614_nl = MUX_s_1_2_2(mux_1613_nl, mux_1612_nl, epsilon_rsci_idat);
  assign mux_1615_nl = MUX_s_1_2_2(mux_1614_nl, or_tmp_210, shift_reg_1_sva_2);
  assign mux_tmp_308 = MUX_s_1_2_2(mux_1620_nl, mux_1615_nl, first_sva);
  assign or_tmp_227 = (~ saved_reg_sva_0) | saved_reg_sva_1 | not_tmp_91;
  assign not_tmp_154 = ~(epsilon_rsci_idat & saved_reg_sva_1 & (count_sva==10'b1111111111));
  assign mux_1626_nl = MUX_s_1_2_2(not_tmp_91, or_tmp_227, epsilon_rsci_idat);
  assign mux_tmp_314 = MUX_s_1_2_2(not_tmp_154, mux_1626_nl, saved_reg_sva_2);
  assign or_tmp_229 = (~(saved_reg_sva_2 & epsilon_rsci_idat & saved_reg_sva_0 &
      (~ saved_reg_sva_1))) | not_tmp_91;
  assign or_tmp_231 = (~ epsilon_rsci_idat) | (~ saved_reg_sva_0) | saved_reg_sva_1
      | not_tmp_91;
  assign mux_1629_nl = MUX_s_1_2_2(not_tmp_154, or_tmp_231, saved_reg_sva_2);
  assign mux_tmp_317 = MUX_s_1_2_2(or_tmp_229, mux_1629_nl, shift_reg_1_sva_0);
  assign mux_tmp_319 = MUX_s_1_2_2(nand_116_cse, or_tmp_100, shift_reg_1_sva_2);
  assign nor_tmp_52 = shift_reg_1_sva_2 & epsilon_rsci_idat;
  assign nand_137_nl = ~(shift_reg_1_sva_0 & shift_reg_1_sva_2 & epsilon_rsci_idat
      & (count_sva==10'b1111111111));
  assign not_tmp_160 = MUX_s_1_2_2(mux_tmp_317, nand_137_nl, first_sva);
  assign mux_1634_nl = MUX_s_1_2_2((~ or_tmp_231), epsilon_rsci_idat, shift_reg_1_sva_2);
  assign mux_1635_nl = MUX_s_1_2_2(nor_tmp_52, mux_1634_nl, saved_reg_sva_2);
  assign mux_1636_nl = MUX_s_1_2_2((~ mux_1635_nl), mux_tmp_314, shift_reg_1_sva_0);
  assign mux_1633_nl = MUX_s_1_2_2((~ nor_tmp_52), mux_tmp_319, shift_reg_1_sva_0);
  assign mux_1637_nl = MUX_s_1_2_2(mux_1636_nl, mux_1633_nl, first_sva);
  assign mux_tmp_326 = MUX_s_1_2_2(not_tmp_160, mux_1637_nl, shift_reg_1_sva_1);
  assign mux_1642_nl = MUX_s_1_2_2(not_tmp_91, or_tmp_227, nor_tmp_52);
  assign mux_tmp_330 = MUX_s_1_2_2(not_tmp_154, mux_1642_nl, saved_reg_sva_2);
  assign and_tmp_12 = shift_reg_1_sva_2 & or_tmp_100;
  assign mux_1648_nl = MUX_s_1_2_2((~ or_tmp_231), or_tmp_100, shift_reg_1_sva_2);
  assign mux_1649_nl = MUX_s_1_2_2(and_tmp_12, mux_1648_nl, saved_reg_sva_2);
  assign mux_1650_nl = MUX_s_1_2_2((~ mux_1649_nl), mux_tmp_330, shift_reg_1_sva_0);
  assign mux_1646_nl = MUX_s_1_2_2(not_tmp_91, mux_tmp_319, saved_reg_sva_2);
  assign mux_1647_nl = MUX_s_1_2_2((~ and_tmp_12), mux_1646_nl, shift_reg_1_sva_0);
  assign mux_1651_nl = MUX_s_1_2_2(mux_1650_nl, mux_1647_nl, first_sva);
  assign mux_tmp_339 = MUX_s_1_2_2(not_tmp_160, mux_1651_nl, shift_reg_1_sva_1);
  assign or_tmp_240 = (~ saved_reg_sva_0) | saved_reg_sva_1 | not_tmp_104;
  assign or_476_nl = (~ saved_reg_sva_1) | saved_reg_sva_2 | (~ and_276_cse);
  assign mux_1658_nl = MUX_s_1_2_2(or_tmp_240, or_476_nl, epsilon_rsci_idat);
  assign mux_1657_nl = MUX_s_1_2_2(not_tmp_104, or_tmp_240, shift_reg_1_sva_1);
  assign or_474_nl = epsilon_rsci_idat | mux_1657_nl;
  assign mux_tmp_346 = MUX_s_1_2_2(mux_1658_nl, or_474_nl, shift_reg_1_sva_0);
  assign or_tmp_245 = first_sva | (~ saved_reg_sva_0) | saved_reg_sva_1 | not_tmp_104;
  assign or_613_nl = first_sva | not_tmp_104;
  assign nand_139_nl = ~(or_tmp_133 & (count_sva==10'b1111111111));
  assign mux_1660_nl = MUX_s_1_2_2(or_613_nl, nand_139_nl, shift_reg_1_sva_2);
  assign mux_1661_nl = MUX_s_1_2_2(mux_1660_nl, or_tmp_245, shift_reg_1_sva_1);
  assign or_tmp_248 = epsilon_rsci_idat | mux_1661_nl;
  assign or_482_cse = (~ shift_reg_1_sva_1) | shift_reg_1_sva_2;
  assign and_tmp_13 = or_482_cse & (first_sva | (~ saved_reg_sva_1) | saved_reg_sva_2
      | (~ and_276_cse));
  assign mux_1662_nl = MUX_s_1_2_2(or_tmp_245, and_tmp_13, epsilon_rsci_idat);
  assign mux_tmp_350 = MUX_s_1_2_2(mux_1662_nl, or_tmp_248, shift_reg_1_sva_0);
  assign nor_195_nl = ~(saved_reg_sva_2 | (~ and_276_cse));
  assign or_488_nl = first_sva | (~ saved_reg_sva_0) | saved_reg_sva_1;
  assign mux_1666_nl = MUX_s_1_2_2(nor_195_nl, and_276_cse, or_488_nl);
  assign mux_1667_nl = MUX_s_1_2_2(mux_1666_nl, or_tmp_245, or_482_cse);
  assign mux_1668_nl = MUX_s_1_2_2(mux_1667_nl, and_tmp_13, epsilon_rsci_idat);
  assign mux_tmp_356 = MUX_s_1_2_2(mux_1668_nl, or_tmp_248, shift_reg_1_sva_0);
  assign mux_tmp_361 = MUX_s_1_2_2(nand_128_cse, or_446_cse, saved_reg_sva_1);
  assign mux_tmp_362 = MUX_s_1_2_2(nand_125_cse, mux_tmp_361, saved_reg_sva_2);
  assign nand_tmp_19 = ~(epsilon_rsci_idat & (~ mux_tmp_362));
  assign not_tmp_175 = ~(shift_reg_1_sva_2 & shift_reg_1_sva_1 & shift_reg_1_sva_0);
  assign mux_1676_nl = MUX_s_1_2_2(nand_128_cse, or_tmp_161, shift_reg_1_sva_1);
  assign mux_1677_nl = MUX_s_1_2_2(nand_125_cse, mux_1676_nl, shift_reg_1_sva_2);
  assign mux_1678_nl = MUX_s_1_2_2(mux_tmp_362, mux_1677_nl, first_sva);
  assign mux_tmp_366 = MUX_s_1_2_2(not_tmp_175, mux_1678_nl, epsilon_rsci_idat);
  assign mux_1685_nl = MUX_s_1_2_2(or_446_cse, and_317_cse, shift_reg_1_sva_0);
  assign mux_1686_nl = MUX_s_1_2_2((~ shift_reg_1_sva_0), mux_1685_nl, saved_reg_sva_1);
  assign mux_1687_nl = MUX_s_1_2_2(mux_tmp_361, mux_1686_nl, shift_reg_1_sva_1);
  assign mux_1688_nl = MUX_s_1_2_2(or_dcpl_65, mux_1687_nl, saved_reg_sva_2);
  assign mux_1689_nl = MUX_s_1_2_2(mux_tmp_362, mux_1688_nl, shift_reg_1_sva_2);
  assign mux_1683_nl = MUX_s_1_2_2(nand_128_cse, mux_1558_cse, shift_reg_1_sva_1);
  assign mux_1684_nl = MUX_s_1_2_2(nand_125_cse, mux_1683_nl, shift_reg_1_sva_2);
  assign mux_1690_nl = MUX_s_1_2_2(mux_1689_nl, mux_1684_nl, first_sva);
  assign mux_tmp_378 = MUX_s_1_2_2(not_tmp_175, mux_1690_nl, epsilon_rsci_idat);
  assign or_tmp_269 = (~ saved_reg_sva_2) | (~ saved_reg_sva_1) | saved_reg_sva_0
      | epsilon_rsci_idat | not_tmp_91;
  assign nor_196_nl = ~(saved_reg_sva_0 | epsilon_rsci_idat | not_tmp_91);
  assign mux_1696_nl = MUX_s_1_2_2(and_294_cse, nor_196_nl, saved_reg_sva_1);
  assign nand_tmp_20 = ~(saved_reg_sva_2 & mux_1696_nl);
  assign or_506_nl = (~ saved_reg_sva_1) | saved_reg_sva_0 | epsilon_rsci_idat |
      not_tmp_91;
  assign mux_tmp_385 = MUX_s_1_2_2((~ and_294_cse), or_506_nl, saved_reg_sva_2);
  assign mux_1699_nl = MUX_s_1_2_2(nand_tmp_20, mux_tmp_385, shift_reg_1_sva_0);
  assign mux_1697_nl = MUX_s_1_2_2(nand_tmp_20, or_tmp_269, shift_reg_1_sva_0);
  assign mux_tmp_387 = MUX_s_1_2_2(mux_1699_nl, mux_1697_nl, shift_reg_1_sva_1);
  assign mux_tmp_390 = MUX_s_1_2_2(nand_tmp_20, or_341_cse, first_sva);
  assign nand_145_nl = ~(shift_reg_1_sva_2 & epsilon_rsci_idat & (count_sva==10'b1111111111));
  assign mux_1706_nl = MUX_s_1_2_2(nand_tmp_20, nand_145_nl, first_sva);
  assign or_510_nl = shift_reg_1_sva_2 | (~ and_294_cse);
  assign mux_1705_nl = MUX_s_1_2_2(mux_tmp_385, or_510_nl, first_sva);
  assign mux_tmp_394 = MUX_s_1_2_2(mux_1706_nl, mux_1705_nl, shift_reg_1_sva_0);
  assign mux_1701_nl = MUX_s_1_2_2(epsilon_rsci_idat, or_tmp_269, shift_reg_1_sva_2);
  assign mux_1702_nl = MUX_s_1_2_2(mux_1701_nl, or_tmp_105, first_sva);
  assign mux_1704_nl = MUX_s_1_2_2(mux_tmp_390, mux_1702_nl, shift_reg_1_sva_0);
  assign mux_tmp_395 = MUX_s_1_2_2(mux_tmp_394, mux_1704_nl, shift_reg_1_sva_1);
  assign mux_1711_nl = MUX_s_1_2_2(and_294_cse, or_tmp_269, shift_reg_1_sva_2);
  assign mux_1712_nl = MUX_s_1_2_2(mux_1711_nl, or_387_cse, first_sva);
  assign mux_1713_nl = MUX_s_1_2_2(mux_tmp_390, mux_1712_nl, shift_reg_1_sva_0);
  assign mux_tmp_401 = MUX_s_1_2_2(mux_tmp_394, mux_1713_nl, shift_reg_1_sva_1);
  assign not_tmp_188 = ~(saved_reg_sva_1 & saved_reg_sva_2 & (count_sva==10'b1111111111));
  assign nor_197_nl = ~((~ saved_reg_sva_0) | first_sva | not_tmp_188);
  assign nor_198_nl = ~(first_sva | not_tmp_188);
  assign or_519_nl = shift_reg_1_sva_2 | (~(first_sva | not_tmp_104));
  assign mux_1720_nl = MUX_s_1_2_2(nor_198_nl, or_519_nl, shift_reg_1_sva_1);
  assign mux_tmp_408 = MUX_s_1_2_2(nor_197_nl, mux_1720_nl, shift_reg_1_sva_0);
  assign and_351_cse = saved_reg_sva_0 & saved_reg_sva_1 & saved_reg_sva_2 & (count_sva==10'b1111111111);
  assign and_352_nl = (shift_reg_1_sva_1 | saved_reg_sva_1) & saved_reg_sva_2 & (count_sva==10'b1111111111);
  assign mux_1719_nl = MUX_s_1_2_2(and_351_cse, and_352_nl, shift_reg_1_sva_0);
  assign mux_1722_nl = MUX_s_1_2_2(mux_tmp_408, mux_1719_nl, or_325_cse);
  assign mux_tmp_410 = MUX_s_1_2_2(mux_tmp_408, mux_1722_nl, or_324_cse);
  assign or_tmp_294 = (~ saved_reg_sva_2) | shift_reg_1_sva_1 | (~ and_276_cse);
  assign nor_tmp_78 = saved_reg_sva_1 & saved_reg_sva_2 & (count_sva==10'b1111111111);
  assign mux_1728_nl = MUX_s_1_2_2((~ nor_tmp_78), or_tmp_294, shift_reg_1_sva_0);
  assign mux_tmp_416 = MUX_s_1_2_2((~ and_351_cse), mux_1728_nl, epsilon_rsci_idat);
  assign nor_tmp_80 = shift_reg_1_sva_2 & shift_reg_1_sva_1 & (count_sva==10'b1111111111);
  assign mux_1734_nl = MUX_s_1_2_2(nor_tmp_78, nor_tmp_80, first_sva);
  assign mux_1731_nl = MUX_s_1_2_2(shift_reg_1_sva_1, or_tmp_93, saved_reg_sva_2);
  assign mux_1732_nl = MUX_s_1_2_2((~ mux_1731_nl), or_tmp_294, shift_reg_1_sva_2);
  assign mux_1730_nl = MUX_s_1_2_2((~ shift_reg_1_sva_1), or_327_cse, shift_reg_1_sva_2);
  assign mux_1733_nl = MUX_s_1_2_2(mux_1732_nl, mux_1730_nl, first_sva);
  assign mux_tmp_422 = MUX_s_1_2_2((~ mux_1734_nl), mux_1733_nl, shift_reg_1_sva_0);
  assign not_tmp_199 = ~(first_sva | (~ and_351_cse));
  assign mux_1736_nl = MUX_s_1_2_2(and_351_cse, nor_tmp_80, first_sva);
  assign mux_1737_nl = MUX_s_1_2_2(not_tmp_199, mux_1736_nl, shift_reg_1_sva_0);
  assign mux_tmp_425 = MUX_s_1_2_2((~ mux_1737_nl), mux_tmp_422, epsilon_rsci_idat);
  assign and_359_nl = saved_reg_sva_0 & saved_reg_sva_1 & saved_reg_sva_2;
  assign mux_1742_nl = MUX_s_1_2_2(not_tmp_88, or_tmp_93, and_359_nl);
  assign mux_1743_nl = MUX_s_1_2_2(mux_1742_nl, and_351_cse, shift_reg_1_sva_2);
  assign and_360_nl = shift_reg_1_sva_1 & (count_sva==10'b1111111111);
  assign mux_1741_nl = MUX_s_1_2_2(not_tmp_88, and_360_nl, shift_reg_1_sva_2);
  assign mux_1744_nl = MUX_s_1_2_2(mux_1743_nl, mux_1741_nl, first_sva);
  assign mux_1745_nl = MUX_s_1_2_2(not_tmp_199, mux_1744_nl, shift_reg_1_sva_0);
  assign mux_tmp_433 = MUX_s_1_2_2((~ mux_1745_nl), mux_tmp_422, epsilon_rsci_idat);
  assign mux_1752_nl = MUX_s_1_2_2(or_dcpl_100, or_tmp_89, first_sva);
  assign mux_1751_nl = MUX_s_1_2_2(or_dcpl_100, or_tmp_89, nor_159_cse);
  assign mux_tmp_440 = MUX_s_1_2_2(mux_1752_nl, mux_1751_nl, or_324_cse);
  assign nand_150_cse = ~(or_324_cse & (skip_sva_1_1_0_1[1]));
  assign or_tmp_306 = ~(nand_150_cse & shift_reg_1_sva_1);
  assign mux_1755_nl = MUX_s_1_2_2(saved_reg_sva_2, shift_reg_1_sva_2, first_sva);
  assign mux_1754_nl = MUX_s_1_2_2(saved_reg_sva_2, shift_reg_1_sva_2, nor_159_cse);
  assign mux_1756_cse = MUX_s_1_2_2(mux_1755_nl, mux_1754_nl, or_324_cse);
  assign mux_tmp_444 = MUX_s_1_2_2(or_tmp_306, mux_1756_cse, shift_reg_1_sva_0);
  assign or_tmp_308 = (~ shift_reg_1_sva_2) | shift_reg_1_sva_1;
  assign or_tmp_309 = shift_reg_1_sva_1 | (~ or_dcpl_100);
  assign or_tmp_310 = ~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_1_3_0_lpi_1_dfm_2_2_0==3'b100)
      & (~ exit_if_4_for_lpi_1_dfm_2));
  assign and_tmp_15 = (skip_sva_1_1_0_1[1]) & or_324_cse;
  assign or_tmp_323 = (~ saved_reg_sva_1) | saved_reg_sva_2;
  assign or_tmp_325 = shift_reg_1_sva_1 | (~ or_tmp_323);
  assign mux_1778_nl = MUX_s_1_2_2(or_tmp_325, shift_reg_1_sva_1, first_sva);
  assign mux_1776_nl = MUX_s_1_2_2(or_tmp_325, shift_reg_1_sva_1, nor_149_cse);
  assign mux_1777_nl = MUX_s_1_2_2((~ mux_1776_nl), or_tmp_323, skip_sva_1_1_0_1[1]);
  assign mux_1779_nl = MUX_s_1_2_2((~ mux_1778_nl), mux_1777_nl, or_324_cse);
  assign mux_1774_nl = MUX_s_1_2_2(or_tmp_323, or_482_cse, first_sva);
  assign mux_1773_nl = MUX_s_1_2_2(or_tmp_323, or_482_cse, nor_159_cse);
  assign mux_1775_nl = MUX_s_1_2_2(mux_1774_nl, mux_1773_nl, or_324_cse);
  assign mux_tmp_467 = MUX_s_1_2_2(mux_1779_nl, mux_1775_nl, shift_reg_1_sva_0);
  assign or_tmp_329 = ~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_1_3_0_lpi_1_dfm_2_2_0==3'b101)
      & (~ exit_if_4_for_lpi_1_dfm_2));
  assign or_tmp_334 = and_tmp_15 | shift_reg_1_sva_1 | shift_reg_1_sva_0;
  assign mux_tmp_479 = MUX_s_1_2_2((~ shift_reg_1_sva_1), shift_reg_1_sva_0, shift_reg_1_sva_2);
  assign mux_tmp_480 = MUX_s_1_2_2((~ saved_reg_sva_1), shift_reg_1_sva_0, saved_reg_sva_2);
  assign or_tmp_336 = ~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_1_3_0_lpi_1_dfm_2_2_0==3'b001)
      & (~ exit_if_4_for_lpi_1_dfm_2));
  assign mux_tmp_485 = MUX_s_1_2_2(or_tmp_336, or_tmp_334, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign nor_205_nl = ~(shift_reg_1_sva_1 | (~ shift_reg_1_sva_0));
  assign mux_tmp_486 = MUX_s_1_2_2(nor_205_nl, shift_reg_1_sva_0, shift_reg_1_sva_2);
  assign nor_206_nl = ~(saved_reg_sva_1 | (~ or_dcpl_26));
  assign mux_tmp_487 = MUX_s_1_2_2(nor_206_nl, shift_reg_1_sva_0, saved_reg_sva_2);
  assign mux_tmp_497 = MUX_s_1_2_2((~ shift_reg_1_sva_0), shift_reg_1_sva_1, shift_reg_1_sva_2);
  assign mux_tmp_498 = MUX_s_1_2_2((~ shift_reg_1_sva_0), saved_reg_sva_1, saved_reg_sva_2);
  assign or_tmp_343 = and_tmp_15 | or_dcpl_65;
  assign or_tmp_346 = nor_87_cse | shift_reg_1_sva_0;
  assign nand_84_nl = ~(saved_reg_sva_1 & or_dcpl_65);
  assign mux_tmp_503 = MUX_s_1_2_2(shift_reg_1_sva_0, nand_84_nl, saved_reg_sva_2);
  assign or_tmp_347 = ~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_1_3_0_lpi_1_dfm_2_2_0==3'b110)
      & (~ exit_if_4_for_lpi_1_dfm_2));
  assign mux_tmp_509 = MUX_s_1_2_2(or_tmp_347, or_tmp_343, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign and_tmp_17 = shift_reg_1_sva_1 & or_tmp_21;
  assign mux_1835_nl = MUX_s_1_2_2(or_tmp_21, or_tmp_308, first_sva);
  assign mux_1834_nl = MUX_s_1_2_2(or_tmp_21, or_tmp_308, nor_159_cse);
  assign mux_1836_nl = MUX_s_1_2_2(mux_1835_nl, mux_1834_nl, or_324_cse);
  assign mux_1832_nl = MUX_s_1_2_2(and_tmp_17, shift_reg_1_sva_1, first_sva);
  assign mux_1830_nl = MUX_s_1_2_2(and_tmp_17, shift_reg_1_sva_1, nor_149_cse);
  assign mux_1831_nl = MUX_s_1_2_2(mux_1830_nl, or_tmp_21, skip_sva_1_1_0_1[1]);
  assign mux_1833_nl = MUX_s_1_2_2(mux_1832_nl, mux_1831_nl, or_324_cse);
  assign mux_tmp_524 = MUX_s_1_2_2(mux_1836_nl, mux_1833_nl, shift_reg_1_sva_0);
  assign or_tmp_356 = and_tmp_15 | shift_reg_1_sva_1;
  assign or_tmp_357 = ~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_1_3_0_lpi_1_dfm_2_2_0==3'b010)
      & (~ exit_if_4_for_lpi_1_dfm_2));
  assign nor_tmp_112 = shift_reg_1_sva_1 & shift_reg_1_sva_0;
  assign mux_tmp_533 = MUX_s_1_2_2(nor_tmp_112, or_dcpl_26, shift_reg_1_sva_2);
  assign mux_tmp_534 = MUX_s_1_2_2(nor_tmp_112, or_tmp_216, saved_reg_sva_2);
  assign mux_1850_nl = MUX_s_1_2_2(mux_tmp_534, mux_tmp_533, first_sva);
  assign mux_1848_nl = MUX_s_1_2_2(mux_tmp_534, mux_tmp_533, nor_149_cse);
  assign and_262_nl = saved_reg_sva_2 & or_tmp_216;
  assign mux_1849_nl = MUX_s_1_2_2(mux_1848_nl, and_262_nl, skip_sva_1_1_0_1[1]);
  assign mux_tmp_538 = MUX_s_1_2_2(mux_1850_nl, mux_1849_nl, or_324_cse);
  assign not_tmp_236 = nand_150_cse & nor_tmp_112;
  assign mux_tmp_546 = MUX_s_1_2_2((~ mux_1756_cse), or_tmp_356, shift_reg_1_sva_0);
  assign nor_tmp_119 = shift_reg_1_sva_2 & shift_reg_1_sva_1;
  assign mux_1861_nl = MUX_s_1_2_2(nor_tmp_5, nor_tmp_119, first_sva);
  assign mux_1860_nl = MUX_s_1_2_2(nor_tmp_5, nor_tmp_119, nor_159_cse);
  assign mux_tmp_549 = MUX_s_1_2_2(mux_1861_nl, mux_1860_nl, or_324_cse);
  assign nand_tmp_28 = ~(shift_reg_1_sva_1 & (~ nor_tmp_5));
  assign or_tmp_370 = ~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_1_3_0_lpi_1_dfm_2_2_0==3'b011)
      & (~ exit_if_4_for_lpi_1_dfm_2));
  assign nor_187_nl = ~(or_dcpl_26 | and_tmp_15);
  assign mux_1770_nl = MUX_s_1_2_2(and_298_cse, nor_187_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign nor_188_nl = ~(or_tmp_209 | and_tmp_15);
  assign mux_1771_nl = MUX_s_1_2_2(mux_1770_nl, nor_188_nl, exitL_exit_approx_sva);
  assign or_548_nl = or_2_tmp | and_298_cse;
  assign mux_1772_ssc = MUX_s_1_2_2(mux_1771_nl, or_548_nl, and_276_cse);
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      is_random_rsci_idat <= 1'b0;
    end
    else if ( ~ or_dcpl_10 ) begin
      is_random_rsci_idat <= (readslicef_14_1_13(if_4_aelse_acc_nl)) & if_4_slc_if_4_acc_1_15_svs_1
          & if_4_for_and_mdf_sva_2 & (~ unequal_tmp_2_2);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      valid_rsci_idat <= 1'b0;
    end
    else if ( ~ or_dcpl_10 ) begin
      valid_rsci_idat <= if_4_for_and_mdf_sva_2 & (~ unequal_tmp_2_2);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      reg_is_random_triosy_obj_ld_cse <= 1'b0;
      exitL_exit_if_4_for_2_lpi_1_dfm_st_1_2 <= 1'b0;
      mux_1304_itm_2 <= 1'b0;
      first_sva <= 1'b1;
      epsilon_triosy_obj_ld <= 1'b0;
      exitL_exit_if_4_for_2_lpi_1_dfm <= 1'b0;
      exitL_exit_approx_sva <= 1'b1;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      mux_1304_itm_1 <= 1'b0;
    end
    else begin
      reg_is_random_triosy_obj_ld_cse <= main_stage_0_3 & exitL_exit_if_4_for_2_lpi_1_dfm_st_1_2;
      exitL_exit_if_4_for_2_lpi_1_dfm_st_1_2 <= exitL_exit_if_4_for_2_lpi_1_dfm;
      mux_1304_itm_2 <= mux_1304_itm_1;
      first_sva <= (first_sva & (~((skip_sva_dfm_1_0_mx0==2'b00) & or_2_tmp))) |
          and_91_tmp_1;
      epsilon_triosy_obj_ld <= ~ and_dcpl_67;
      exitL_exit_if_4_for_2_lpi_1_dfm <= exitL_exit_if_4_for_2_lpi_1_dfm_1;
      exitL_exit_approx_sva <= exitL_exit_if_4_for_2_lpi_1_dfm_1;
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
      mux_1304_itm_1 <= MUX_s_1_2_2(if_4_for_if_4_for_or_4_nl, or_2_tmp, nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_4_aelse_not_itm_1 <= 13'b0000000000000;
    end
    else if ( (asn_sft_lpi_1_dfm_st_1==10'b1111111111) & main_stage_0_2 & if_4_for_and_mdf_sva_st_1
        & if_4_acc_1_itm_15_1 & mux_1304_itm_1 ) begin
      if_4_aelse_not_itm_1 <= ~ (if_4_acc_psp_sva_1[14:2]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_4_slc_if_4_acc_1_15_svs_1 <= 1'b0;
      if_4_for_and_mdf_sva_2 <= 1'b0;
      unequal_tmp_2_2 <= 1'b0;
    end
    else if ( and_dcpl_24 ) begin
      if_4_slc_if_4_acc_1_15_svs_1 <= MUX_s_1_2_2(if_4_acc_1_itm_15_1, if_4_slc_if_4_acc_1_15_svs,
          or_40_nl);
      if_4_for_and_mdf_sva_2 <= if_4_for_and_mdf_sva_st_1;
      unequal_tmp_2_2 <= unequal_tmp_2_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      sum1_1_lpi_1_dfm_1 <= 24'b000000000000000000000000;
    end
    else if ( MUX_s_1_2_2(and_275_nl, and_276_cse, or_2_tmp) ) begin
      sum1_1_lpi_1_dfm_1 <= MUX_v_24_2_2(24'b000000000000000000000000, sum1_1_lpi_1_dfm_2_mx0,
          if_4_for_if_4_for_if_4_for_not_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      ln_land_251_lpi_1_dfm_1 <= 1'b0;
      ln_land_252_lpi_1_dfm_1 <= 1'b0;
      ln_ln_mux1h_118_psp_1_12 <= 1'b0;
      ln_and_248_ssc_1 <= 1'b0;
      ln_if_253_acc_cse_11_sva_1 <= 1'b0;
      ln_ln_mux1h_118_psp_1_11 <= 1'b0;
      ln_ln_mux1h_118_psp_1_10 <= 1'b0;
      ln_and_407_ssc_1 <= 1'b0;
      ln_and_244_ssc_1 <= 1'b0;
      ln_and_379_ssc_1 <= 1'b0;
      ln_and_240_ssc_1 <= 1'b0;
      ln_and_377_ssc_1 <= 1'b0;
      ln_and_242_ssc_1 <= 1'b0;
      ln_and_427_itm_1 <= 1'b0;
      ln_ln_mux1h_118_psp_1_8 <= 1'b0;
      ln_ln_mux1h_118_psp_1_7 <= 1'b0;
      ln_ln_mux1h_118_psp_1_6 <= 1'b0;
      ln_ln_mux1h_118_psp_1_5 <= 1'b0;
      ln_ln_mux1h_118_psp_1_4 <= 1'b0;
      ln_ln_mux1h_118_psp_1_3 <= 1'b0;
      ln_ln_mux1h_118_psp_1_2 <= 1'b0;
      ln_ln_mux1h_118_psp_1_1 <= 1'b0;
      ln_ln_mux1h_118_psp_1_0 <= 1'b0;
      operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1 <= 14'b00000000000000;
    end
    else if ( and_dcpl_49 ) begin
      ln_land_251_lpi_1_dfm_1 <= ln_land_251_lpi_1_dfm_1_1;
      ln_land_252_lpi_1_dfm_1 <= ln_land_252_lpi_1_dfm_1_1;
      ln_ln_mux1h_118_psp_1_12 <= (~(ln_land_141_lpi_1_dfm_1 | ln_land_142_lpi_1_dfm_1))
          & ln_nor_3_cse_1 & (~(ln_and_140_ssc_1 | ln_land_146_lpi_1_dfm_1 | ln_land_147_lpi_1_dfm_1
          | ln_land_148_lpi_1_dfm_1 | ln_land_149_lpi_1_dfm_1 | ln_land_150_lpi_1_dfm_1
          | ln_land_151_lpi_1_dfm_1 | ln_land_152_lpi_1_dfm_1 | ln_land_153_lpi_1_dfm_1
          | ln_land_154_lpi_1_dfm_1 | ln_land_155_lpi_1_dfm_1 | ln_land_156_lpi_1_dfm_1
          | ln_land_157_lpi_1_dfm_1 | ln_land_158_lpi_1_dfm_1 | ln_land_159_lpi_1_dfm_1
          | ln_land_160_lpi_1_dfm_1 | ln_land_161_lpi_1_dfm_1 | ln_land_162_lpi_1_dfm_1
          | ln_land_163_lpi_1_dfm_1 | ln_land_164_lpi_1_dfm_1 | ln_land_165_lpi_1_dfm_1
          | ln_land_166_lpi_1_dfm_1 | ln_land_167_lpi_1_dfm_1 | ln_land_168_lpi_1_dfm_1
          | ln_land_169_lpi_1_dfm_1 | ln_land_170_lpi_1_dfm_1 | ln_land_171_lpi_1_dfm_1
          | ln_land_172_lpi_1_dfm_1 | ln_land_173_lpi_1_dfm_1 | ln_land_174_lpi_1_dfm_1
          | ln_land_175_lpi_1_dfm_1 | ln_land_176_lpi_1_dfm_1 | ln_land_177_lpi_1_dfm_1
          | ln_land_178_lpi_1_dfm_1 | ln_land_179_lpi_1_dfm_1 | ln_land_180_lpi_1_dfm_1
          | ln_land_181_lpi_1_dfm_1 | ln_land_182_lpi_1_dfm_1 | ln_land_183_lpi_1_dfm_1
          | ln_land_184_lpi_1_dfm_1 | ln_land_185_lpi_1_dfm_1 | ln_land_186_lpi_1_dfm_1
          | ln_land_187_lpi_1_dfm_1 | ln_land_188_lpi_1_dfm_1 | ln_land_189_lpi_1_dfm_1
          | ln_land_190_lpi_1_dfm_1 | ln_land_191_lpi_1_dfm_1 | ln_land_192_lpi_1_dfm_1
          | ln_land_193_lpi_1_dfm_1 | ln_land_194_lpi_1_dfm_1 | ln_land_195_lpi_1_dfm_1
          | ln_land_196_lpi_1_dfm_1 | ln_land_197_lpi_1_dfm_1 | ln_land_198_lpi_1_dfm_1
          | ln_land_199_lpi_1_dfm_1 | ln_land_200_lpi_1_dfm_1 | ln_land_201_lpi_1_dfm_1
          | ln_land_202_lpi_1_dfm_1 | ln_land_203_lpi_1_dfm_1 | ln_land_204_lpi_1_dfm_1
          | ln_land_205_lpi_1_dfm_1 | ln_land_206_lpi_1_dfm_1 | ln_land_207_lpi_1_dfm_1
          | ln_land_208_lpi_1_dfm_1 | ln_land_209_lpi_1_dfm_1 | ln_land_210_lpi_1_dfm_1
          | ln_land_211_lpi_1_dfm_1 | ln_land_212_lpi_1_dfm_1 | ln_land_213_lpi_1_dfm_1
          | ln_land_214_lpi_1_dfm_1 | ln_land_215_lpi_1_dfm_1 | ln_land_216_lpi_1_dfm_1
          | ln_land_217_lpi_1_dfm_1 | ln_land_218_lpi_1_dfm_1 | ln_land_219_lpi_1_dfm_1
          | ln_land_220_lpi_1_dfm_1 | ln_land_221_lpi_1_dfm_1 | ln_land_222_lpi_1_dfm_1
          | ln_land_223_lpi_1_dfm_1 | ln_land_224_lpi_1_dfm_1 | ln_land_225_lpi_1_dfm_1
          | ln_land_226_lpi_1_dfm_1 | ln_land_227_lpi_1_dfm_1 | ln_land_228_lpi_1_dfm_1
          | ln_land_229_lpi_1_dfm_1 | ln_land_230_lpi_1_dfm_1 | ln_land_231_lpi_1_dfm_1
          | ln_land_232_lpi_1_dfm_1 | ln_land_233_lpi_1_dfm_1 | ln_land_234_lpi_1_dfm_1
          | ln_land_235_lpi_1_dfm_1 | ln_land_236_lpi_1_dfm_1 | ln_land_237_lpi_1_dfm_1
          | ln_land_238_lpi_1_dfm_1 | ln_land_239_lpi_1_dfm_1 | ln_land_240_lpi_1_dfm_1
          | ln_land_241_lpi_1_dfm_1 | ln_land_242_lpi_1_dfm_1 | ln_land_243_lpi_1_dfm_1
          | ln_land_244_lpi_1_dfm_1));
      ln_and_248_ssc_1 <= ln_if_252_acc_itm_12_1 & (~ ln_if_253_acc_itm_11_1);
      ln_if_253_acc_cse_11_sva_1 <= ln_if_253_acc_itm_11_1;
      ln_ln_mux1h_118_psp_1_11 <= ((((~(ln_land_51_lpi_1_dfm_1 | ln_land_52_lpi_1_dfm_1))
          & (~(ln_and_48_ssc_1 | ln_land_54_lpi_1_dfm_1 | ln_land_55_lpi_1_dfm_1
          | ln_land_56_lpi_1_dfm_1 | ln_land_57_lpi_1_dfm_1 | ln_land_58_lpi_1_dfm_1
          | ln_land_59_lpi_1_dfm_1 | ln_land_60_lpi_1_dfm_1 | ln_land_61_lpi_1_dfm_1
          | ln_land_62_lpi_1_dfm_1 | ln_land_63_lpi_1_dfm_1 | ln_land_64_lpi_1_dfm_1
          | ln_land_65_lpi_1_dfm_1 | ln_land_66_lpi_1_dfm_1 | ln_land_67_lpi_1_dfm_1
          | ln_land_68_lpi_1_dfm_1 | ln_land_69_lpi_1_dfm_1 | ln_land_70_lpi_1_dfm_1
          | ln_land_71_lpi_1_dfm_1 | ln_land_72_lpi_1_dfm_1 | ln_land_73_lpi_1_dfm_1
          | ln_land_74_lpi_1_dfm_1 | ln_land_75_lpi_1_dfm_1 | ln_land_76_lpi_1_dfm_1
          | ln_land_77_lpi_1_dfm_1 | ln_land_78_lpi_1_dfm_1 | ln_land_79_lpi_1_dfm_1
          | ln_land_80_lpi_1_dfm_1 | ln_land_81_lpi_1_dfm_1 | ln_land_82_lpi_1_dfm_1
          | ln_land_83_lpi_1_dfm_1 | ln_land_84_lpi_1_dfm_1 | ln_land_85_lpi_1_dfm_1
          | ln_land_86_lpi_1_dfm_1 | ln_land_87_lpi_1_dfm_1 | ln_land_88_lpi_1_dfm_1
          | ln_land_89_lpi_1_dfm_1 | ln_land_90_lpi_1_dfm_1 | ln_land_91_lpi_1_dfm_1
          | ln_land_92_lpi_1_dfm_1 | ln_land_93_lpi_1_dfm_1 | ln_land_94_lpi_1_dfm_1
          | ln_land_95_lpi_1_dfm_1 | ln_land_96_lpi_1_dfm_1 | ln_land_97_lpi_1_dfm_1
          | ln_land_98_lpi_1_dfm_1 | ln_land_99_lpi_1_dfm_1 | ln_land_100_lpi_1_dfm_1
          | ln_land_101_lpi_1_dfm_1 | ln_land_102_lpi_1_dfm_1 | ln_land_103_lpi_1_dfm_1
          | ln_land_104_lpi_1_dfm_1 | ln_land_105_lpi_1_dfm_1 | ln_land_106_lpi_1_dfm_1
          | ln_land_107_lpi_1_dfm_1 | ln_land_108_lpi_1_dfm_1 | ln_land_109_lpi_1_dfm_1
          | ln_land_110_lpi_1_dfm_1 | ln_land_111_lpi_1_dfm_1 | ln_land_112_lpi_1_dfm_1
          | ln_land_113_lpi_1_dfm_1 | ln_land_114_lpi_1_dfm_1 | ln_land_115_lpi_1_dfm_1
          | ln_land_116_lpi_1_dfm_1 | ln_land_117_lpi_1_dfm_1 | ln_land_118_lpi_1_dfm_1
          | ln_land_119_lpi_1_dfm_1 | ln_land_120_lpi_1_dfm_1 | ln_land_121_lpi_1_dfm_1
          | ln_land_122_lpi_1_dfm_1 | ln_land_123_lpi_1_dfm_1 | ln_land_124_lpi_1_dfm_1
          | ln_land_125_lpi_1_dfm_1 | ln_land_126_lpi_1_dfm_1 | ln_land_127_lpi_1_dfm_1
          | ln_land_128_lpi_1_dfm_1 | ln_land_129_lpi_1_dfm_1 | ln_land_130_lpi_1_dfm_1
          | ln_land_131_lpi_1_dfm_1 | ln_land_132_lpi_1_dfm_1 | ln_land_133_lpi_1_dfm_1
          | ln_land_134_lpi_1_dfm_1 | ln_land_135_lpi_1_dfm_1 | ln_land_136_lpi_1_dfm_1
          | ln_land_137_lpi_1_dfm_1 | ln_land_138_lpi_1_dfm_1 | ln_land_139_lpi_1_dfm_1
          | ln_land_140_lpi_1_dfm_1))) | ln_land_141_lpi_1_dfm_1 | ln_land_142_lpi_1_dfm_1
          | ln_and_138_ssc_1 | ln_land_144_lpi_1_dfm_1) & ln_and_368_m1c_1) | ln_and_140_ssc_1
          | ln_land_146_lpi_1_dfm_1 | ln_land_147_lpi_1_dfm_1 | ln_land_148_lpi_1_dfm_1
          | ln_land_149_lpi_1_dfm_1 | ln_land_150_lpi_1_dfm_1 | ln_land_151_lpi_1_dfm_1
          | ln_land_152_lpi_1_dfm_1 | ln_land_153_lpi_1_dfm_1 | ln_land_154_lpi_1_dfm_1
          | ln_land_155_lpi_1_dfm_1 | ln_land_156_lpi_1_dfm_1 | ln_land_157_lpi_1_dfm_1
          | ln_land_158_lpi_1_dfm_1 | ln_land_159_lpi_1_dfm_1 | ln_land_160_lpi_1_dfm_1
          | ln_land_161_lpi_1_dfm_1 | ln_land_162_lpi_1_dfm_1 | ln_land_163_lpi_1_dfm_1
          | ln_land_164_lpi_1_dfm_1 | ln_land_165_lpi_1_dfm_1 | ln_land_166_lpi_1_dfm_1
          | ln_land_167_lpi_1_dfm_1 | ln_land_168_lpi_1_dfm_1 | ln_land_169_lpi_1_dfm_1
          | ln_land_170_lpi_1_dfm_1 | ln_land_171_lpi_1_dfm_1 | ln_land_172_lpi_1_dfm_1
          | ln_land_173_lpi_1_dfm_1 | ln_land_174_lpi_1_dfm_1 | ln_land_175_lpi_1_dfm_1
          | ln_land_176_lpi_1_dfm_1 | ln_land_177_lpi_1_dfm_1 | ln_land_178_lpi_1_dfm_1
          | ln_land_179_lpi_1_dfm_1 | ln_land_180_lpi_1_dfm_1 | ln_land_181_lpi_1_dfm_1
          | ln_land_182_lpi_1_dfm_1 | ln_land_183_lpi_1_dfm_1 | ln_land_184_lpi_1_dfm_1
          | ln_land_185_lpi_1_dfm_1 | ln_land_186_lpi_1_dfm_1 | ln_land_187_lpi_1_dfm_1
          | ln_land_188_lpi_1_dfm_1 | ln_land_189_lpi_1_dfm_1 | ln_land_190_lpi_1_dfm_1
          | ln_land_191_lpi_1_dfm_1 | ln_land_192_lpi_1_dfm_1 | ln_land_193_lpi_1_dfm_1
          | ln_land_194_lpi_1_dfm_1 | ln_land_195_lpi_1_dfm_1 | ln_land_196_lpi_1_dfm_1
          | ln_land_197_lpi_1_dfm_1 | ln_land_198_lpi_1_dfm_1 | ln_land_199_lpi_1_dfm_1
          | ln_land_200_lpi_1_dfm_1 | ln_land_201_lpi_1_dfm_1 | ln_land_202_lpi_1_dfm_1
          | ln_land_203_lpi_1_dfm_1 | ln_land_204_lpi_1_dfm_1 | ln_land_205_lpi_1_dfm_1
          | ln_land_206_lpi_1_dfm_1 | ln_land_207_lpi_1_dfm_1 | ln_land_208_lpi_1_dfm_1
          | ln_land_209_lpi_1_dfm_1 | ln_land_210_lpi_1_dfm_1 | ln_land_211_lpi_1_dfm_1
          | ln_land_212_lpi_1_dfm_1 | ln_land_213_lpi_1_dfm_1 | ln_land_214_lpi_1_dfm_1
          | ln_land_215_lpi_1_dfm_1 | ln_land_216_lpi_1_dfm_1 | ln_land_217_lpi_1_dfm_1
          | ln_land_218_lpi_1_dfm_1 | ln_land_219_lpi_1_dfm_1 | ln_land_220_lpi_1_dfm_1
          | ln_land_221_lpi_1_dfm_1 | ln_land_222_lpi_1_dfm_1 | ln_land_223_lpi_1_dfm_1
          | ln_land_224_lpi_1_dfm_1 | ln_land_225_lpi_1_dfm_1 | ln_land_226_lpi_1_dfm_1
          | ln_land_227_lpi_1_dfm_1 | ln_land_228_lpi_1_dfm_1;
      ln_ln_mux1h_118_psp_1_10 <= (((((~(ln_land_6_lpi_1_dfm_1 | ln_and_4_ssc_1 |
          ln_land_8_lpi_1_dfm_1 | ln_land_9_lpi_1_dfm_1 | ln_land_10_lpi_1_dfm_1
          | ln_land_11_lpi_1_dfm_1 | ln_land_12_lpi_1_dfm_1 | ln_land_13_lpi_1_dfm_1
          | ln_land_14_lpi_1_dfm_1 | ln_land_15_lpi_1_dfm_1 | ln_land_16_lpi_1_dfm_1
          | ln_land_17_lpi_1_dfm_1 | ln_land_18_lpi_1_dfm_1 | ln_land_19_lpi_1_dfm_1
          | ln_land_20_lpi_1_dfm_1 | ln_land_21_lpi_1_dfm_1 | ln_land_22_lpi_1_dfm_1
          | ln_land_23_lpi_1_dfm_1 | ln_land_24_lpi_1_dfm_1 | ln_land_25_lpi_1_dfm_1
          | ln_land_26_lpi_1_dfm_1 | ln_land_27_lpi_1_dfm_1 | ln_land_28_lpi_1_dfm_1
          | ln_land_29_lpi_1_dfm_1 | ln_land_30_lpi_1_dfm_1 | ln_land_31_lpi_1_dfm_1
          | ln_land_32_lpi_1_dfm_1 | ln_land_33_lpi_1_dfm_1 | ln_land_34_lpi_1_dfm_1
          | ln_land_35_lpi_1_dfm_1 | ln_land_36_lpi_1_dfm_1 | ln_land_37_lpi_1_dfm_1
          | ln_land_38_lpi_1_dfm_1 | ln_land_39_lpi_1_dfm_1 | ln_land_40_lpi_1_dfm_1
          | ln_land_41_lpi_1_dfm_1 | ln_land_42_lpi_1_dfm_1 | ln_land_43_lpi_1_dfm_1
          | ln_land_44_lpi_1_dfm_1 | ln_land_45_lpi_1_dfm_1 | ln_land_46_lpi_1_dfm_1
          | ln_land_47_lpi_1_dfm_1 | ln_land_48_lpi_1_dfm_1 | ln_land_49_lpi_1_dfm_1
          | ln_if_50_ln_if_50_and_seb_1)) | ln_land_51_lpi_1_dfm_1 | ln_land_52_lpi_1_dfm_1)
          & (~(ln_land_98_lpi_1_dfm_1 | ln_land_99_lpi_1_dfm_1 | ln_land_100_lpi_1_dfm_1
          | ln_land_101_lpi_1_dfm_1 | ln_land_102_lpi_1_dfm_1 | ln_land_103_lpi_1_dfm_1
          | ln_land_104_lpi_1_dfm_1 | ln_land_105_lpi_1_dfm_1 | ln_land_106_lpi_1_dfm_1
          | ln_land_107_lpi_1_dfm_1 | ln_land_108_lpi_1_dfm_1 | ln_land_109_lpi_1_dfm_1
          | ln_land_110_lpi_1_dfm_1 | ln_land_111_lpi_1_dfm_1 | ln_land_112_lpi_1_dfm_1
          | ln_land_113_lpi_1_dfm_1 | ln_land_114_lpi_1_dfm_1 | ln_land_115_lpi_1_dfm_1
          | ln_land_116_lpi_1_dfm_1 | ln_land_117_lpi_1_dfm_1 | ln_land_118_lpi_1_dfm_1
          | ln_land_119_lpi_1_dfm_1 | ln_land_120_lpi_1_dfm_1 | ln_land_121_lpi_1_dfm_1
          | ln_land_122_lpi_1_dfm_1 | ln_land_123_lpi_1_dfm_1 | ln_land_124_lpi_1_dfm_1
          | ln_land_125_lpi_1_dfm_1 | ln_land_126_lpi_1_dfm_1 | ln_land_127_lpi_1_dfm_1
          | ln_land_128_lpi_1_dfm_1 | ln_land_129_lpi_1_dfm_1 | ln_land_130_lpi_1_dfm_1
          | ln_land_131_lpi_1_dfm_1 | ln_land_132_lpi_1_dfm_1 | ln_land_133_lpi_1_dfm_1
          | ln_land_134_lpi_1_dfm_1 | ln_land_135_lpi_1_dfm_1 | ln_land_136_lpi_1_dfm_1
          | ln_land_137_lpi_1_dfm_1 | ln_land_138_lpi_1_dfm_1 | ln_land_139_lpi_1_dfm_1
          | ln_land_140_lpi_1_dfm_1))) | ln_and_48_ssc_1 | ln_land_54_lpi_1_dfm_1
          | ln_land_55_lpi_1_dfm_1 | ln_land_56_lpi_1_dfm_1 | ln_land_57_lpi_1_dfm_1
          | ln_land_58_lpi_1_dfm_1 | ln_land_59_lpi_1_dfm_1 | ln_land_60_lpi_1_dfm_1
          | ln_land_61_lpi_1_dfm_1 | ln_land_62_lpi_1_dfm_1 | ln_land_63_lpi_1_dfm_1
          | ln_land_64_lpi_1_dfm_1 | ln_land_65_lpi_1_dfm_1 | ln_land_66_lpi_1_dfm_1
          | ln_land_67_lpi_1_dfm_1 | ln_land_68_lpi_1_dfm_1 | ln_land_69_lpi_1_dfm_1
          | ln_land_70_lpi_1_dfm_1 | ln_land_71_lpi_1_dfm_1 | ln_land_72_lpi_1_dfm_1
          | ln_land_73_lpi_1_dfm_1 | ln_land_74_lpi_1_dfm_1 | ln_land_75_lpi_1_dfm_1
          | ln_land_76_lpi_1_dfm_1 | ln_land_77_lpi_1_dfm_1 | ln_land_78_lpi_1_dfm_1
          | ln_land_79_lpi_1_dfm_1 | ln_land_80_lpi_1_dfm_1 | ln_land_81_lpi_1_dfm_1
          | ln_land_82_lpi_1_dfm_1 | ln_land_83_lpi_1_dfm_1 | ln_land_84_lpi_1_dfm_1
          | ln_land_85_lpi_1_dfm_1 | ln_land_86_lpi_1_dfm_1 | ln_land_87_lpi_1_dfm_1
          | ln_land_88_lpi_1_dfm_1 | ln_land_89_lpi_1_dfm_1 | ln_land_90_lpi_1_dfm_1
          | ln_land_91_lpi_1_dfm_1 | ln_land_92_lpi_1_dfm_1 | ln_land_93_lpi_1_dfm_1
          | ln_land_94_lpi_1_dfm_1 | ln_land_95_lpi_1_dfm_1 | ln_land_96_lpi_1_dfm_1
          | ln_land_97_lpi_1_dfm_1 | ln_land_141_lpi_1_dfm_1 | ln_land_142_lpi_1_dfm_1
          | ln_and_138_ssc_1 | ln_land_144_lpi_1_dfm_1) & (~(ln_land_195_lpi_1_dfm_1
          | ln_land_196_lpi_1_dfm_1 | ln_land_197_lpi_1_dfm_1 | ln_land_198_lpi_1_dfm_1
          | ln_land_199_lpi_1_dfm_1 | ln_land_200_lpi_1_dfm_1 | ln_land_201_lpi_1_dfm_1
          | ln_land_202_lpi_1_dfm_1 | ln_land_203_lpi_1_dfm_1 | ln_land_204_lpi_1_dfm_1
          | ln_land_205_lpi_1_dfm_1 | ln_land_206_lpi_1_dfm_1 | ln_land_207_lpi_1_dfm_1
          | ln_land_208_lpi_1_dfm_1 | ln_land_209_lpi_1_dfm_1 | ln_land_210_lpi_1_dfm_1
          | ln_land_211_lpi_1_dfm_1 | ln_land_212_lpi_1_dfm_1 | ln_land_213_lpi_1_dfm_1
          | ln_land_214_lpi_1_dfm_1 | ln_land_215_lpi_1_dfm_1 | ln_land_216_lpi_1_dfm_1
          | ln_land_217_lpi_1_dfm_1 | ln_land_218_lpi_1_dfm_1 | ln_land_219_lpi_1_dfm_1
          | ln_land_220_lpi_1_dfm_1 | ln_land_221_lpi_1_dfm_1 | ln_land_222_lpi_1_dfm_1
          | ln_land_223_lpi_1_dfm_1 | ln_land_224_lpi_1_dfm_1 | ln_land_225_lpi_1_dfm_1
          | ln_land_226_lpi_1_dfm_1 | ln_land_227_lpi_1_dfm_1 | ln_land_228_lpi_1_dfm_1)))
          | ln_and_140_ssc_1 | ln_land_146_lpi_1_dfm_1 | ln_land_147_lpi_1_dfm_1
          | ln_land_148_lpi_1_dfm_1 | ln_land_149_lpi_1_dfm_1 | ln_land_150_lpi_1_dfm_1
          | ln_land_151_lpi_1_dfm_1 | ln_land_152_lpi_1_dfm_1 | ln_land_153_lpi_1_dfm_1
          | ln_land_154_lpi_1_dfm_1 | ln_land_155_lpi_1_dfm_1 | ln_land_156_lpi_1_dfm_1
          | ln_land_157_lpi_1_dfm_1 | ln_land_158_lpi_1_dfm_1 | ln_land_159_lpi_1_dfm_1
          | ln_land_160_lpi_1_dfm_1 | ln_land_161_lpi_1_dfm_1 | ln_land_162_lpi_1_dfm_1
          | ln_land_163_lpi_1_dfm_1 | ln_land_164_lpi_1_dfm_1 | ln_land_165_lpi_1_dfm_1
          | ln_land_166_lpi_1_dfm_1 | ln_land_167_lpi_1_dfm_1 | ln_land_168_lpi_1_dfm_1
          | ln_land_169_lpi_1_dfm_1 | ln_land_170_lpi_1_dfm_1 | ln_land_171_lpi_1_dfm_1
          | ln_land_172_lpi_1_dfm_1 | ln_land_173_lpi_1_dfm_1 | ln_land_174_lpi_1_dfm_1
          | ln_land_175_lpi_1_dfm_1 | ln_land_176_lpi_1_dfm_1 | ln_land_177_lpi_1_dfm_1
          | ln_land_178_lpi_1_dfm_1 | ln_land_179_lpi_1_dfm_1 | ln_land_180_lpi_1_dfm_1
          | ln_land_181_lpi_1_dfm_1 | ln_land_182_lpi_1_dfm_1 | ln_land_183_lpi_1_dfm_1
          | ln_land_184_lpi_1_dfm_1 | ln_land_185_lpi_1_dfm_1 | ln_land_186_lpi_1_dfm_1
          | ln_land_187_lpi_1_dfm_1 | ln_land_188_lpi_1_dfm_1 | ln_land_189_lpi_1_dfm_1
          | ln_land_190_lpi_1_dfm_1 | ln_land_191_lpi_1_dfm_1 | ln_land_192_lpi_1_dfm_1
          | ln_land_193_lpi_1_dfm_1 | ln_land_194_lpi_1_dfm_1 | ln_land_229_lpi_1_dfm_1
          | ln_land_230_lpi_1_dfm_1 | ln_land_231_lpi_1_dfm_1 | ln_land_232_lpi_1_dfm_1
          | ln_land_233_lpi_1_dfm_1 | ln_land_234_lpi_1_dfm_1 | ln_land_235_lpi_1_dfm_1
          | ln_land_236_lpi_1_dfm_1 | ln_land_237_lpi_1_dfm_1 | ln_land_238_lpi_1_dfm_1
          | ln_land_239_lpi_1_dfm_1 | ln_land_240_lpi_1_dfm_1 | ln_land_241_lpi_1_dfm_1
          | ln_land_242_lpi_1_dfm_1 | ln_land_243_lpi_1_dfm_1 | ln_land_244_lpi_1_dfm_1;
      ln_and_407_ssc_1 <= ln_land_248_lpi_1_dfm_1;
      ln_and_244_ssc_1 <= ln_land_249_lpi_1_dfm_1;
      ln_and_379_ssc_1 <= ln_land_250_lpi_1_dfm_1;
      ln_and_240_ssc_1 <= ln_and_240_ssc_1_1;
      ln_and_377_ssc_1 <= ln_land_246_lpi_1_dfm_1;
      ln_and_242_ssc_1 <= ln_land_247_lpi_1_dfm_1;
      ln_and_427_itm_1 <= ((((((~(ln_nor_33_cse_1 | ln_land_17_lpi_1_dfm_1 | ln_land_18_lpi_1_dfm_1
          | ln_land_19_lpi_1_dfm_1 | ln_land_20_lpi_1_dfm_1 | ln_land_21_lpi_1_dfm_1
          | ln_land_22_lpi_1_dfm_1 | ln_land_23_lpi_1_dfm_1 | ln_land_24_lpi_1_dfm_1
          | ln_land_25_lpi_1_dfm_1 | ln_land_26_lpi_1_dfm_1 | ln_land_27_lpi_1_dfm_1
          | ln_land_28_lpi_1_dfm_1 | ln_land_29_lpi_1_dfm_1 | ln_land_30_lpi_1_dfm_1
          | ln_land_31_lpi_1_dfm_1 | ln_land_32_lpi_1_dfm_1 | ln_land_33_lpi_1_dfm_1
          | ln_land_34_lpi_1_dfm_1 | ln_land_35_lpi_1_dfm_1 | ln_land_36_lpi_1_dfm_1
          | ln_land_37_lpi_1_dfm_1 | ln_land_38_lpi_1_dfm_1 | ln_land_39_lpi_1_dfm_1
          | ln_land_40_lpi_1_dfm_1 | ln_land_41_lpi_1_dfm_1 | ln_land_42_lpi_1_dfm_1
          | ln_land_43_lpi_1_dfm_1 | ln_land_44_lpi_1_dfm_1 | ln_land_45_lpi_1_dfm_1
          | ln_land_46_lpi_1_dfm_1 | ln_land_47_lpi_1_dfm_1 | ln_land_48_lpi_1_dfm_1
          | ln_land_49_lpi_1_dfm_1 | ln_if_50_ln_if_50_and_seb_1)) | ln_land_51_lpi_1_dfm_1
          | ln_land_52_lpi_1_dfm_1) & (~(ln_land_77_lpi_1_dfm_1 | ln_land_78_lpi_1_dfm_1
          | ln_land_79_lpi_1_dfm_1 | ln_land_80_lpi_1_dfm_1 | ln_land_81_lpi_1_dfm_1
          | ln_land_82_lpi_1_dfm_1 | ln_land_83_lpi_1_dfm_1 | ln_land_84_lpi_1_dfm_1
          | ln_land_85_lpi_1_dfm_1 | ln_land_86_lpi_1_dfm_1 | ln_land_87_lpi_1_dfm_1
          | ln_land_88_lpi_1_dfm_1 | ln_land_89_lpi_1_dfm_1 | ln_land_90_lpi_1_dfm_1
          | ln_land_91_lpi_1_dfm_1 | ln_land_92_lpi_1_dfm_1 | ln_land_93_lpi_1_dfm_1
          | ln_land_94_lpi_1_dfm_1 | ln_land_95_lpi_1_dfm_1 | ln_land_96_lpi_1_dfm_1
          | ln_land_97_lpi_1_dfm_1 | ln_land_114_lpi_1_dfm_1 | ln_land_115_lpi_1_dfm_1
          | ln_land_116_lpi_1_dfm_1 | ln_land_117_lpi_1_dfm_1 | ln_land_118_lpi_1_dfm_1
          | ln_land_119_lpi_1_dfm_1 | ln_land_120_lpi_1_dfm_1 | ln_land_121_lpi_1_dfm_1
          | ln_land_122_lpi_1_dfm_1 | ln_land_123_lpi_1_dfm_1 | ln_land_124_lpi_1_dfm_1
          | ln_land_125_lpi_1_dfm_1 | ln_land_126_lpi_1_dfm_1 | ln_land_127_lpi_1_dfm_1
          | ln_land_128_lpi_1_dfm_1 | ln_land_129_lpi_1_dfm_1 | ln_land_130_lpi_1_dfm_1
          | ln_land_131_lpi_1_dfm_1 | ln_land_132_lpi_1_dfm_1 | ln_land_133_lpi_1_dfm_1
          | ln_land_134_lpi_1_dfm_1 | ln_land_135_lpi_1_dfm_1 | ln_land_136_lpi_1_dfm_1
          | ln_land_137_lpi_1_dfm_1 | ln_land_138_lpi_1_dfm_1 | ln_land_139_lpi_1_dfm_1
          | ln_land_140_lpi_1_dfm_1))) | ln_and_48_ssc_1 | ln_land_54_lpi_1_dfm_1
          | ln_land_55_lpi_1_dfm_1 | ln_land_56_lpi_1_dfm_1 | ln_land_57_lpi_1_dfm_1
          | ln_land_58_lpi_1_dfm_1 | ln_land_59_lpi_1_dfm_1 | ln_land_60_lpi_1_dfm_1
          | ln_land_61_lpi_1_dfm_1 | ln_land_62_lpi_1_dfm_1 | ln_land_63_lpi_1_dfm_1
          | ln_land_64_lpi_1_dfm_1 | ln_land_65_lpi_1_dfm_1 | ln_land_66_lpi_1_dfm_1
          | ln_land_67_lpi_1_dfm_1 | ln_land_68_lpi_1_dfm_1 | ln_land_69_lpi_1_dfm_1
          | ln_land_70_lpi_1_dfm_1 | ln_land_71_lpi_1_dfm_1 | ln_land_72_lpi_1_dfm_1
          | ln_land_73_lpi_1_dfm_1 | ln_land_74_lpi_1_dfm_1 | ln_land_75_lpi_1_dfm_1
          | ln_land_76_lpi_1_dfm_1 | ln_land_98_lpi_1_dfm_1 | ln_land_99_lpi_1_dfm_1
          | ln_land_100_lpi_1_dfm_1 | ln_land_101_lpi_1_dfm_1 | ln_land_102_lpi_1_dfm_1
          | ln_land_103_lpi_1_dfm_1 | ln_land_104_lpi_1_dfm_1 | ln_land_105_lpi_1_dfm_1
          | ln_land_106_lpi_1_dfm_1 | ln_land_107_lpi_1_dfm_1 | ln_land_108_lpi_1_dfm_1
          | ln_land_109_lpi_1_dfm_1 | ln_land_110_lpi_1_dfm_1 | ln_land_111_lpi_1_dfm_1
          | ln_land_112_lpi_1_dfm_1 | ln_land_113_lpi_1_dfm_1 | ln_land_141_lpi_1_dfm_1
          | ln_land_142_lpi_1_dfm_1 | ln_and_138_ssc_1 | ln_land_144_lpi_1_dfm_1)
          & (~(ln_land_172_lpi_1_dfm_1 | ln_land_173_lpi_1_dfm_1 | ln_land_174_lpi_1_dfm_1
          | ln_land_175_lpi_1_dfm_1 | ln_land_176_lpi_1_dfm_1 | ln_land_177_lpi_1_dfm_1
          | ln_land_178_lpi_1_dfm_1 | ln_land_179_lpi_1_dfm_1 | ln_land_180_lpi_1_dfm_1
          | ln_land_181_lpi_1_dfm_1 | ln_land_182_lpi_1_dfm_1 | ln_land_183_lpi_1_dfm_1
          | ln_land_184_lpi_1_dfm_1 | ln_land_185_lpi_1_dfm_1 | ln_land_186_lpi_1_dfm_1
          | ln_land_187_lpi_1_dfm_1 | ln_land_188_lpi_1_dfm_1 | ln_land_189_lpi_1_dfm_1
          | ln_land_190_lpi_1_dfm_1 | ln_land_191_lpi_1_dfm_1 | ln_land_192_lpi_1_dfm_1
          | ln_land_193_lpi_1_dfm_1 | ln_land_194_lpi_1_dfm_1 | ln_land_214_lpi_1_dfm_1
          | ln_land_215_lpi_1_dfm_1 | ln_land_216_lpi_1_dfm_1 | ln_land_217_lpi_1_dfm_1
          | ln_land_218_lpi_1_dfm_1 | ln_land_219_lpi_1_dfm_1 | ln_land_220_lpi_1_dfm_1
          | ln_land_221_lpi_1_dfm_1 | ln_land_222_lpi_1_dfm_1 | ln_land_223_lpi_1_dfm_1
          | ln_land_224_lpi_1_dfm_1 | ln_land_225_lpi_1_dfm_1 | ln_land_226_lpi_1_dfm_1
          | ln_land_227_lpi_1_dfm_1 | ln_land_228_lpi_1_dfm_1 | ln_land_240_lpi_1_dfm_1
          | ln_land_241_lpi_1_dfm_1 | ln_land_242_lpi_1_dfm_1 | ln_land_243_lpi_1_dfm_1
          | ln_land_244_lpi_1_dfm_1))) | ln_and_140_ssc_1 | ln_land_146_lpi_1_dfm_1
          | ln_land_147_lpi_1_dfm_1 | ln_land_148_lpi_1_dfm_1 | ln_land_149_lpi_1_dfm_1
          | ln_land_150_lpi_1_dfm_1 | ln_land_151_lpi_1_dfm_1 | ln_land_152_lpi_1_dfm_1
          | ln_land_153_lpi_1_dfm_1 | ln_land_154_lpi_1_dfm_1 | ln_land_155_lpi_1_dfm_1
          | ln_land_156_lpi_1_dfm_1 | ln_land_157_lpi_1_dfm_1 | ln_land_158_lpi_1_dfm_1
          | ln_land_159_lpi_1_dfm_1 | ln_land_160_lpi_1_dfm_1 | ln_land_161_lpi_1_dfm_1
          | ln_land_162_lpi_1_dfm_1 | ln_land_163_lpi_1_dfm_1 | ln_land_164_lpi_1_dfm_1
          | ln_land_165_lpi_1_dfm_1 | ln_land_166_lpi_1_dfm_1 | ln_land_167_lpi_1_dfm_1
          | ln_land_168_lpi_1_dfm_1 | ln_land_169_lpi_1_dfm_1 | ln_land_170_lpi_1_dfm_1
          | ln_land_171_lpi_1_dfm_1 | ln_land_195_lpi_1_dfm_1 | ln_land_196_lpi_1_dfm_1
          | ln_land_197_lpi_1_dfm_1 | ln_land_198_lpi_1_dfm_1 | ln_land_199_lpi_1_dfm_1
          | ln_land_200_lpi_1_dfm_1 | ln_land_201_lpi_1_dfm_1 | ln_land_202_lpi_1_dfm_1
          | ln_land_203_lpi_1_dfm_1 | ln_land_204_lpi_1_dfm_1 | ln_land_205_lpi_1_dfm_1
          | ln_land_206_lpi_1_dfm_1 | ln_land_207_lpi_1_dfm_1 | ln_land_208_lpi_1_dfm_1
          | ln_land_209_lpi_1_dfm_1 | ln_land_210_lpi_1_dfm_1 | ln_land_211_lpi_1_dfm_1
          | ln_land_212_lpi_1_dfm_1 | ln_land_213_lpi_1_dfm_1 | ln_land_229_lpi_1_dfm_1
          | ln_land_230_lpi_1_dfm_1 | ln_land_231_lpi_1_dfm_1 | ln_land_232_lpi_1_dfm_1
          | ln_land_233_lpi_1_dfm_1 | ln_land_234_lpi_1_dfm_1 | ln_land_235_lpi_1_dfm_1
          | ln_land_236_lpi_1_dfm_1 | ln_land_237_lpi_1_dfm_1 | ln_land_238_lpi_1_dfm_1
          | ln_land_239_lpi_1_dfm_1) & (~(ln_and_240_ssc_1_1 | ln_land_246_lpi_1_dfm_1
          | ln_land_247_lpi_1_dfm_1 | ln_land_249_lpi_1_dfm_1 | ln_land_250_lpi_1_dfm_1
          | ln_land_252_lpi_1_dfm_1_1));
      ln_ln_mux1h_118_psp_1_8 <= (((((~(((~((~(ln_nor_5_cse_1 | ln_and_2_ssc_1))
          | ln_land_6_lpi_1_dfm_1)) & (~(ln_land_17_lpi_1_dfm_1 | ln_land_18_lpi_1_dfm_1
          | ln_land_19_lpi_1_dfm_1 | ln_land_20_lpi_1_dfm_1 | ln_land_21_lpi_1_dfm_1
          | ln_land_22_lpi_1_dfm_1 | ln_land_23_lpi_1_dfm_1 | ln_land_24_lpi_1_dfm_1
          | ln_land_25_lpi_1_dfm_1 | ln_land_26_lpi_1_dfm_1 | ln_land_27_lpi_1_dfm_1
          | ln_land_28_lpi_1_dfm_1 | ln_land_29_lpi_1_dfm_1 | ln_land_30_lpi_1_dfm_1
          | ln_land_31_lpi_1_dfm_1 | ln_land_32_lpi_1_dfm_1 | ln_land_33_lpi_1_dfm_1
          | ln_land_34_lpi_1_dfm_1))) | ln_and_4_ssc_1 | ln_land_8_lpi_1_dfm_1 |
          ln_land_9_lpi_1_dfm_1 | ln_land_10_lpi_1_dfm_1 | ln_land_11_lpi_1_dfm_1
          | ln_land_12_lpi_1_dfm_1 | ln_land_13_lpi_1_dfm_1 | ln_land_14_lpi_1_dfm_1
          | ln_land_15_lpi_1_dfm_1 | ln_land_16_lpi_1_dfm_1 | ln_land_35_lpi_1_dfm_1
          | ln_land_36_lpi_1_dfm_1 | ln_land_37_lpi_1_dfm_1 | ln_land_38_lpi_1_dfm_1
          | ln_land_39_lpi_1_dfm_1 | ln_land_40_lpi_1_dfm_1 | ln_land_41_lpi_1_dfm_1
          | ln_land_42_lpi_1_dfm_1 | ln_land_43_lpi_1_dfm_1 | ln_land_44_lpi_1_dfm_1
          | ln_land_45_lpi_1_dfm_1 | ln_land_46_lpi_1_dfm_1 | ln_land_47_lpi_1_dfm_1
          | ln_land_48_lpi_1_dfm_1 | ln_land_49_lpi_1_dfm_1 | ln_if_50_ln_if_50_and_seb_1))
          | ln_land_51_lpi_1_dfm_1 | ln_land_52_lpi_1_dfm_1) & (~(ln_land_65_lpi_1_dfm_1
          | ln_land_66_lpi_1_dfm_1 | ln_land_67_lpi_1_dfm_1 | ln_land_68_lpi_1_dfm_1
          | ln_land_69_lpi_1_dfm_1 | ln_land_70_lpi_1_dfm_1 | ln_land_71_lpi_1_dfm_1
          | ln_land_72_lpi_1_dfm_1 | ln_land_73_lpi_1_dfm_1 | ln_land_74_lpi_1_dfm_1
          | ln_land_75_lpi_1_dfm_1 | ln_land_76_lpi_1_dfm_1 | ln_land_88_lpi_1_dfm_1
          | ln_land_89_lpi_1_dfm_1 | ln_land_90_lpi_1_dfm_1 | ln_land_91_lpi_1_dfm_1
          | ln_land_92_lpi_1_dfm_1 | ln_land_93_lpi_1_dfm_1 | ln_land_94_lpi_1_dfm_1
          | ln_land_95_lpi_1_dfm_1 | ln_land_96_lpi_1_dfm_1 | ln_land_97_lpi_1_dfm_1
          | ln_land_106_lpi_1_dfm_1 | ln_land_107_lpi_1_dfm_1 | ln_land_108_lpi_1_dfm_1
          | ln_land_109_lpi_1_dfm_1 | ln_land_110_lpi_1_dfm_1 | ln_land_111_lpi_1_dfm_1
          | ln_land_112_lpi_1_dfm_1 | ln_land_113_lpi_1_dfm_1 | ln_land_122_lpi_1_dfm_1
          | ln_land_123_lpi_1_dfm_1 | ln_land_124_lpi_1_dfm_1 | ln_land_125_lpi_1_dfm_1
          | ln_land_126_lpi_1_dfm_1 | ln_land_127_lpi_1_dfm_1 | ln_land_128_lpi_1_dfm_1
          | ln_land_129_lpi_1_dfm_1 | ln_land_130_lpi_1_dfm_1 | ln_land_131_lpi_1_dfm_1
          | ln_land_132_lpi_1_dfm_1 | ln_land_133_lpi_1_dfm_1 | ln_land_134_lpi_1_dfm_1
          | ln_land_135_lpi_1_dfm_1 | ln_land_136_lpi_1_dfm_1 | ln_land_137_lpi_1_dfm_1
          | ln_land_138_lpi_1_dfm_1 | ln_land_139_lpi_1_dfm_1 | ln_land_140_lpi_1_dfm_1)))
          | ln_and_48_ssc_1 | ln_land_54_lpi_1_dfm_1 | ln_land_55_lpi_1_dfm_1 | ln_land_56_lpi_1_dfm_1
          | ln_land_57_lpi_1_dfm_1 | ln_land_58_lpi_1_dfm_1 | ln_land_59_lpi_1_dfm_1
          | ln_land_60_lpi_1_dfm_1 | ln_land_61_lpi_1_dfm_1 | ln_land_62_lpi_1_dfm_1
          | ln_land_63_lpi_1_dfm_1 | ln_land_64_lpi_1_dfm_1 | ln_land_77_lpi_1_dfm_1
          | ln_land_78_lpi_1_dfm_1 | ln_land_79_lpi_1_dfm_1 | ln_land_80_lpi_1_dfm_1
          | ln_land_81_lpi_1_dfm_1 | ln_land_82_lpi_1_dfm_1 | ln_land_83_lpi_1_dfm_1
          | ln_land_84_lpi_1_dfm_1 | ln_land_85_lpi_1_dfm_1 | ln_land_86_lpi_1_dfm_1
          | ln_land_87_lpi_1_dfm_1 | ln_land_98_lpi_1_dfm_1 | ln_land_99_lpi_1_dfm_1
          | ln_land_100_lpi_1_dfm_1 | ln_land_101_lpi_1_dfm_1 | ln_land_102_lpi_1_dfm_1
          | ln_land_103_lpi_1_dfm_1 | ln_land_104_lpi_1_dfm_1 | ln_land_105_lpi_1_dfm_1
          | ln_land_114_lpi_1_dfm_1 | ln_land_115_lpi_1_dfm_1 | ln_land_116_lpi_1_dfm_1
          | ln_land_117_lpi_1_dfm_1 | ln_land_118_lpi_1_dfm_1 | ln_land_119_lpi_1_dfm_1
          | ln_land_120_lpi_1_dfm_1 | ln_land_121_lpi_1_dfm_1 | ln_land_141_lpi_1_dfm_1
          | ln_land_142_lpi_1_dfm_1 | ln_and_138_ssc_1 | ln_land_144_lpi_1_dfm_1)
          & (~(ln_land_157_lpi_1_dfm_1 | ln_land_158_lpi_1_dfm_1 | ln_land_159_lpi_1_dfm_1
          | ln_land_160_lpi_1_dfm_1 | ln_land_161_lpi_1_dfm_1 | ln_land_162_lpi_1_dfm_1
          | ln_land_163_lpi_1_dfm_1 | ln_land_164_lpi_1_dfm_1 | ln_land_165_lpi_1_dfm_1
          | ln_land_166_lpi_1_dfm_1 | ln_land_167_lpi_1_dfm_1 | ln_land_168_lpi_1_dfm_1
          | ln_land_169_lpi_1_dfm_1 | ln_land_170_lpi_1_dfm_1 | ln_land_171_lpi_1_dfm_1
          | ln_land_184_lpi_1_dfm_1 | ln_land_185_lpi_1_dfm_1 | ln_land_186_lpi_1_dfm_1
          | ln_land_187_lpi_1_dfm_1 | ln_land_188_lpi_1_dfm_1 | ln_land_189_lpi_1_dfm_1
          | ln_land_190_lpi_1_dfm_1 | ln_land_191_lpi_1_dfm_1 | ln_land_192_lpi_1_dfm_1
          | ln_land_193_lpi_1_dfm_1 | ln_land_194_lpi_1_dfm_1 | ln_land_205_lpi_1_dfm_1
          | ln_land_206_lpi_1_dfm_1 | ln_land_207_lpi_1_dfm_1 | ln_land_208_lpi_1_dfm_1
          | ln_land_209_lpi_1_dfm_1 | ln_land_210_lpi_1_dfm_1 | ln_land_211_lpi_1_dfm_1
          | ln_land_212_lpi_1_dfm_1 | ln_land_213_lpi_1_dfm_1 | ln_land_222_lpi_1_dfm_1
          | ln_land_223_lpi_1_dfm_1 | ln_land_224_lpi_1_dfm_1 | ln_land_225_lpi_1_dfm_1
          | ln_land_226_lpi_1_dfm_1 | ln_land_227_lpi_1_dfm_1 | ln_land_228_lpi_1_dfm_1
          | ln_land_235_lpi_1_dfm_1 | ln_land_236_lpi_1_dfm_1 | ln_land_237_lpi_1_dfm_1
          | ln_land_238_lpi_1_dfm_1 | ln_land_239_lpi_1_dfm_1 | ln_land_244_lpi_1_dfm_1)))
          | ln_and_140_ssc_1 | ln_land_146_lpi_1_dfm_1 | ln_land_147_lpi_1_dfm_1
          | ln_land_148_lpi_1_dfm_1 | ln_land_149_lpi_1_dfm_1 | ln_land_150_lpi_1_dfm_1
          | ln_land_151_lpi_1_dfm_1 | ln_land_152_lpi_1_dfm_1 | ln_land_153_lpi_1_dfm_1
          | ln_land_154_lpi_1_dfm_1 | ln_land_155_lpi_1_dfm_1 | ln_land_156_lpi_1_dfm_1
          | ln_land_172_lpi_1_dfm_1 | ln_land_173_lpi_1_dfm_1 | ln_land_174_lpi_1_dfm_1
          | ln_land_175_lpi_1_dfm_1 | ln_land_176_lpi_1_dfm_1 | ln_land_177_lpi_1_dfm_1
          | ln_land_178_lpi_1_dfm_1 | ln_land_179_lpi_1_dfm_1 | ln_land_180_lpi_1_dfm_1
          | ln_land_181_lpi_1_dfm_1 | ln_land_182_lpi_1_dfm_1 | ln_land_183_lpi_1_dfm_1
          | ln_land_195_lpi_1_dfm_1 | ln_land_196_lpi_1_dfm_1 | ln_land_197_lpi_1_dfm_1
          | ln_land_198_lpi_1_dfm_1 | ln_land_199_lpi_1_dfm_1 | ln_land_200_lpi_1_dfm_1
          | ln_land_201_lpi_1_dfm_1 | ln_land_202_lpi_1_dfm_1 | ln_land_203_lpi_1_dfm_1
          | ln_land_204_lpi_1_dfm_1 | ln_land_214_lpi_1_dfm_1 | ln_land_215_lpi_1_dfm_1
          | ln_land_216_lpi_1_dfm_1 | ln_land_217_lpi_1_dfm_1 | ln_land_218_lpi_1_dfm_1
          | ln_land_219_lpi_1_dfm_1 | ln_land_220_lpi_1_dfm_1 | ln_land_221_lpi_1_dfm_1
          | ln_land_229_lpi_1_dfm_1 | ln_land_230_lpi_1_dfm_1 | ln_land_231_lpi_1_dfm_1
          | ln_land_232_lpi_1_dfm_1 | ln_land_233_lpi_1_dfm_1 | ln_land_234_lpi_1_dfm_1
          | ln_land_240_lpi_1_dfm_1 | ln_land_241_lpi_1_dfm_1 | ln_land_242_lpi_1_dfm_1
          | ln_land_243_lpi_1_dfm_1;
      ln_ln_mux1h_118_psp_1_7 <= (((((~(((~(ln_ln_ln_nor_8_cse_1 & ln_nor_1_cse_1))
          & (~(ln_land_17_lpi_1_dfm_1 | ln_land_18_lpi_1_dfm_1 | ln_land_19_lpi_1_dfm_1
          | ln_land_20_lpi_1_dfm_1 | ln_land_21_lpi_1_dfm_1 | ln_land_22_lpi_1_dfm_1
          | ln_land_23_lpi_1_dfm_1 | ln_land_24_lpi_1_dfm_1 | ln_land_25_lpi_1_dfm_1
          | ln_land_35_lpi_1_dfm_1 | ln_land_36_lpi_1_dfm_1 | ln_land_37_lpi_1_dfm_1
          | ln_land_38_lpi_1_dfm_1 | ln_land_39_lpi_1_dfm_1 | ln_land_40_lpi_1_dfm_1
          | ln_land_41_lpi_1_dfm_1 | ln_land_42_lpi_1_dfm_1))) | ln_and_4_ssc_1 |
          ln_land_8_lpi_1_dfm_1 | ln_land_9_lpi_1_dfm_1 | ln_land_10_lpi_1_dfm_1
          | ln_land_11_lpi_1_dfm_1 | ln_land_12_lpi_1_dfm_1 | ln_land_13_lpi_1_dfm_1
          | ln_land_14_lpi_1_dfm_1 | ln_land_15_lpi_1_dfm_1 | ln_land_16_lpi_1_dfm_1
          | ln_land_26_lpi_1_dfm_1 | ln_land_27_lpi_1_dfm_1 | ln_land_28_lpi_1_dfm_1
          | ln_land_29_lpi_1_dfm_1 | ln_land_30_lpi_1_dfm_1 | ln_land_31_lpi_1_dfm_1
          | ln_land_32_lpi_1_dfm_1 | ln_land_33_lpi_1_dfm_1 | ln_land_34_lpi_1_dfm_1
          | ln_land_43_lpi_1_dfm_1 | ln_land_44_lpi_1_dfm_1 | ln_land_45_lpi_1_dfm_1
          | ln_land_46_lpi_1_dfm_1 | ln_land_47_lpi_1_dfm_1 | ln_land_48_lpi_1_dfm_1
          | ln_land_49_lpi_1_dfm_1 | ln_if_50_ln_if_50_and_seb_1)) | ln_land_51_lpi_1_dfm_1
          | ln_land_52_lpi_1_dfm_1) & (~(ln_land_58_lpi_1_dfm_1 | ln_land_59_lpi_1_dfm_1
          | ln_land_60_lpi_1_dfm_1 | ln_land_61_lpi_1_dfm_1 | ln_land_62_lpi_1_dfm_1
          | ln_land_63_lpi_1_dfm_1 | ln_land_64_lpi_1_dfm_1 | ln_land_71_lpi_1_dfm_1
          | ln_land_72_lpi_1_dfm_1 | ln_land_73_lpi_1_dfm_1 | ln_land_74_lpi_1_dfm_1
          | ln_land_75_lpi_1_dfm_1 | ln_land_76_lpi_1_dfm_1 | ln_land_83_lpi_1_dfm_1
          | ln_land_84_lpi_1_dfm_1 | ln_land_85_lpi_1_dfm_1 | ln_land_86_lpi_1_dfm_1
          | ln_land_87_lpi_1_dfm_1 | ln_land_93_lpi_1_dfm_1 | ln_land_94_lpi_1_dfm_1
          | ln_land_95_lpi_1_dfm_1 | ln_land_96_lpi_1_dfm_1 | ln_land_97_lpi_1_dfm_1
          | ln_land_102_lpi_1_dfm_1 | ln_land_103_lpi_1_dfm_1 | ln_land_104_lpi_1_dfm_1
          | ln_land_105_lpi_1_dfm_1 | ln_land_110_lpi_1_dfm_1 | ln_land_111_lpi_1_dfm_1
          | ln_land_112_lpi_1_dfm_1 | ln_land_113_lpi_1_dfm_1 | ln_land_117_lpi_1_dfm_1
          | ln_land_118_lpi_1_dfm_1 | ln_land_119_lpi_1_dfm_1 | ln_land_120_lpi_1_dfm_1
          | ln_land_121_lpi_1_dfm_1 | ln_land_132_lpi_1_dfm_1 | ln_land_133_lpi_1_dfm_1
          | ln_land_134_lpi_1_dfm_1 | ln_land_135_lpi_1_dfm_1 | ln_land_136_lpi_1_dfm_1
          | ln_land_137_lpi_1_dfm_1 | ln_land_138_lpi_1_dfm_1 | ln_land_139_lpi_1_dfm_1
          | ln_land_140_lpi_1_dfm_1))) | ln_and_48_ssc_1 | ln_land_54_lpi_1_dfm_1
          | ln_land_55_lpi_1_dfm_1 | ln_land_56_lpi_1_dfm_1 | ln_land_57_lpi_1_dfm_1
          | ln_land_65_lpi_1_dfm_1 | ln_land_66_lpi_1_dfm_1 | ln_land_67_lpi_1_dfm_1
          | ln_land_68_lpi_1_dfm_1 | ln_land_69_lpi_1_dfm_1 | ln_land_70_lpi_1_dfm_1
          | ln_land_77_lpi_1_dfm_1 | ln_land_78_lpi_1_dfm_1 | ln_land_79_lpi_1_dfm_1
          | ln_land_80_lpi_1_dfm_1 | ln_land_81_lpi_1_dfm_1 | ln_land_82_lpi_1_dfm_1
          | ln_land_88_lpi_1_dfm_1 | ln_land_89_lpi_1_dfm_1 | ln_land_90_lpi_1_dfm_1
          | ln_land_91_lpi_1_dfm_1 | ln_land_92_lpi_1_dfm_1 | ln_land_98_lpi_1_dfm_1
          | ln_land_99_lpi_1_dfm_1 | ln_land_100_lpi_1_dfm_1 | ln_land_101_lpi_1_dfm_1
          | ln_land_106_lpi_1_dfm_1 | ln_land_107_lpi_1_dfm_1 | ln_land_108_lpi_1_dfm_1
          | ln_land_109_lpi_1_dfm_1 | ln_land_114_lpi_1_dfm_1 | ln_land_115_lpi_1_dfm_1
          | ln_land_116_lpi_1_dfm_1 | ln_land_122_lpi_1_dfm_1 | ln_land_123_lpi_1_dfm_1
          | ln_land_124_lpi_1_dfm_1 | ln_land_125_lpi_1_dfm_1 | ln_land_126_lpi_1_dfm_1
          | ln_land_127_lpi_1_dfm_1 | ln_land_128_lpi_1_dfm_1 | ln_land_129_lpi_1_dfm_1
          | ln_land_130_lpi_1_dfm_1 | ln_land_131_lpi_1_dfm_1 | ln_land_141_lpi_1_dfm_1
          | ln_land_142_lpi_1_dfm_1 | ln_and_138_ssc_1 | ln_land_144_lpi_1_dfm_1)
          & (~(ln_land_149_lpi_1_dfm_1 | ln_land_150_lpi_1_dfm_1 | ln_land_151_lpi_1_dfm_1
          | ln_land_152_lpi_1_dfm_1 | ln_land_153_lpi_1_dfm_1 | ln_land_154_lpi_1_dfm_1
          | ln_land_155_lpi_1_dfm_1 | ln_land_156_lpi_1_dfm_1 | ln_land_165_lpi_1_dfm_1
          | ln_land_166_lpi_1_dfm_1 | ln_land_167_lpi_1_dfm_1 | ln_land_168_lpi_1_dfm_1
          | ln_land_169_lpi_1_dfm_1 | ln_land_170_lpi_1_dfm_1 | ln_land_171_lpi_1_dfm_1
          | ln_land_178_lpi_1_dfm_1 | ln_land_179_lpi_1_dfm_1 | ln_land_180_lpi_1_dfm_1
          | ln_land_181_lpi_1_dfm_1 | ln_land_182_lpi_1_dfm_1 | ln_land_183_lpi_1_dfm_1
          | ln_land_190_lpi_1_dfm_1 | ln_land_191_lpi_1_dfm_1 | ln_land_192_lpi_1_dfm_1
          | ln_land_193_lpi_1_dfm_1 | ln_land_194_lpi_1_dfm_1 | ln_land_201_lpi_1_dfm_1
          | ln_land_202_lpi_1_dfm_1 | ln_land_203_lpi_1_dfm_1 | ln_land_204_lpi_1_dfm_1
          | ln_land_210_lpi_1_dfm_1 | ln_land_211_lpi_1_dfm_1 | ln_land_212_lpi_1_dfm_1
          | ln_land_213_lpi_1_dfm_1 | ln_land_218_lpi_1_dfm_1 | ln_land_219_lpi_1_dfm_1
          | ln_land_220_lpi_1_dfm_1 | ln_land_221_lpi_1_dfm_1 | ln_land_225_lpi_1_dfm_1
          | ln_land_226_lpi_1_dfm_1 | ln_land_227_lpi_1_dfm_1 | ln_land_228_lpi_1_dfm_1
          | ln_land_232_lpi_1_dfm_1 | ln_land_233_lpi_1_dfm_1 | ln_land_234_lpi_1_dfm_1
          | ln_land_237_lpi_1_dfm_1 | ln_land_238_lpi_1_dfm_1 | ln_land_239_lpi_1_dfm_1
          | ln_land_242_lpi_1_dfm_1 | ln_land_243_lpi_1_dfm_1))) | ln_and_140_ssc_1
          | ln_land_146_lpi_1_dfm_1 | ln_land_147_lpi_1_dfm_1 | ln_land_148_lpi_1_dfm_1
          | ln_land_157_lpi_1_dfm_1 | ln_land_158_lpi_1_dfm_1 | ln_land_159_lpi_1_dfm_1
          | ln_land_160_lpi_1_dfm_1 | ln_land_161_lpi_1_dfm_1 | ln_land_162_lpi_1_dfm_1
          | ln_land_163_lpi_1_dfm_1 | ln_land_164_lpi_1_dfm_1 | ln_land_172_lpi_1_dfm_1
          | ln_land_173_lpi_1_dfm_1 | ln_land_174_lpi_1_dfm_1 | ln_land_175_lpi_1_dfm_1
          | ln_land_176_lpi_1_dfm_1 | ln_land_177_lpi_1_dfm_1 | ln_land_184_lpi_1_dfm_1
          | ln_land_185_lpi_1_dfm_1 | ln_land_186_lpi_1_dfm_1 | ln_land_187_lpi_1_dfm_1
          | ln_land_188_lpi_1_dfm_1 | ln_land_189_lpi_1_dfm_1 | ln_land_195_lpi_1_dfm_1
          | ln_land_196_lpi_1_dfm_1 | ln_land_197_lpi_1_dfm_1 | ln_land_198_lpi_1_dfm_1
          | ln_land_199_lpi_1_dfm_1 | ln_land_200_lpi_1_dfm_1 | ln_land_205_lpi_1_dfm_1
          | ln_land_206_lpi_1_dfm_1 | ln_land_207_lpi_1_dfm_1 | ln_land_208_lpi_1_dfm_1
          | ln_land_209_lpi_1_dfm_1 | ln_land_214_lpi_1_dfm_1 | ln_land_215_lpi_1_dfm_1
          | ln_land_216_lpi_1_dfm_1 | ln_land_217_lpi_1_dfm_1 | ln_land_222_lpi_1_dfm_1
          | ln_land_223_lpi_1_dfm_1 | ln_land_224_lpi_1_dfm_1 | ln_land_229_lpi_1_dfm_1
          | ln_land_230_lpi_1_dfm_1 | ln_land_231_lpi_1_dfm_1 | ln_land_235_lpi_1_dfm_1
          | ln_land_236_lpi_1_dfm_1 | ln_land_240_lpi_1_dfm_1 | ln_land_241_lpi_1_dfm_1
          | ln_land_244_lpi_1_dfm_1;
      ln_ln_mux1h_118_psp_1_6 <= (((((~(ln_nor_33_cse_1 | ln_land_12_lpi_1_dfm_1
          | ln_land_13_lpi_1_dfm_1 | ln_land_14_lpi_1_dfm_1 | ln_land_15_lpi_1_dfm_1
          | ln_land_16_lpi_1_dfm_1 | ln_land_21_lpi_1_dfm_1 | ln_land_22_lpi_1_dfm_1
          | ln_land_23_lpi_1_dfm_1 | ln_land_24_lpi_1_dfm_1 | ln_land_25_lpi_1_dfm_1
          | ln_land_30_lpi_1_dfm_1 | ln_land_31_lpi_1_dfm_1 | ln_land_32_lpi_1_dfm_1
          | ln_land_33_lpi_1_dfm_1 | ln_land_34_lpi_1_dfm_1 | ln_land_39_lpi_1_dfm_1
          | ln_land_40_lpi_1_dfm_1 | ln_land_41_lpi_1_dfm_1 | ln_land_42_lpi_1_dfm_1
          | ln_land_47_lpi_1_dfm_1 | ln_land_48_lpi_1_dfm_1 | ln_land_49_lpi_1_dfm_1
          | ln_if_50_ln_if_50_and_seb_1)) | ln_land_51_lpi_1_dfm_1 | ln_land_52_lpi_1_dfm_1)
          & (~(ln_land_54_lpi_1_dfm_1 | ln_land_55_lpi_1_dfm_1 | ln_land_56_lpi_1_dfm_1
          | ln_land_57_lpi_1_dfm_1 | ln_land_61_lpi_1_dfm_1 | ln_land_62_lpi_1_dfm_1
          | ln_land_63_lpi_1_dfm_1 | ln_land_64_lpi_1_dfm_1 | ln_land_68_lpi_1_dfm_1
          | ln_land_69_lpi_1_dfm_1 | ln_land_70_lpi_1_dfm_1 | ln_land_74_lpi_1_dfm_1
          | ln_land_75_lpi_1_dfm_1 | ln_land_76_lpi_1_dfm_1 | ln_land_80_lpi_1_dfm_1
          | ln_land_81_lpi_1_dfm_1 | ln_land_82_lpi_1_dfm_1 | ln_land_85_lpi_1_dfm_1
          | ln_land_86_lpi_1_dfm_1 | ln_land_87_lpi_1_dfm_1 | ln_land_91_lpi_1_dfm_1
          | ln_land_92_lpi_1_dfm_1 | ln_land_95_lpi_1_dfm_1 | ln_land_96_lpi_1_dfm_1
          | ln_land_97_lpi_1_dfm_1 | ln_land_100_lpi_1_dfm_1 | ln_land_101_lpi_1_dfm_1
          | ln_land_104_lpi_1_dfm_1 | ln_land_105_lpi_1_dfm_1 | ln_land_108_lpi_1_dfm_1
          | ln_land_109_lpi_1_dfm_1 | ln_land_112_lpi_1_dfm_1 | ln_land_113_lpi_1_dfm_1
          | ln_land_116_lpi_1_dfm_1 | ln_land_119_lpi_1_dfm_1 | ln_land_120_lpi_1_dfm_1
          | ln_land_121_lpi_1_dfm_1 | ln_land_127_lpi_1_dfm_1 | ln_land_128_lpi_1_dfm_1
          | ln_land_129_lpi_1_dfm_1 | ln_land_130_lpi_1_dfm_1 | ln_land_131_lpi_1_dfm_1
          | ln_land_137_lpi_1_dfm_1 | ln_land_138_lpi_1_dfm_1 | ln_land_139_lpi_1_dfm_1
          | ln_land_140_lpi_1_dfm_1))) | ln_and_48_ssc_1 | ln_land_58_lpi_1_dfm_1
          | ln_land_59_lpi_1_dfm_1 | ln_land_60_lpi_1_dfm_1 | ln_land_65_lpi_1_dfm_1
          | ln_land_66_lpi_1_dfm_1 | ln_land_67_lpi_1_dfm_1 | ln_land_71_lpi_1_dfm_1
          | ln_land_72_lpi_1_dfm_1 | ln_land_73_lpi_1_dfm_1 | ln_land_77_lpi_1_dfm_1
          | ln_land_78_lpi_1_dfm_1 | ln_land_79_lpi_1_dfm_1 | ln_land_83_lpi_1_dfm_1
          | ln_land_84_lpi_1_dfm_1 | ln_land_88_lpi_1_dfm_1 | ln_land_89_lpi_1_dfm_1
          | ln_land_90_lpi_1_dfm_1 | ln_land_93_lpi_1_dfm_1 | ln_land_94_lpi_1_dfm_1
          | ln_land_98_lpi_1_dfm_1 | ln_land_99_lpi_1_dfm_1 | ln_land_102_lpi_1_dfm_1
          | ln_land_103_lpi_1_dfm_1 | ln_land_106_lpi_1_dfm_1 | ln_land_107_lpi_1_dfm_1
          | ln_land_110_lpi_1_dfm_1 | ln_land_111_lpi_1_dfm_1 | ln_land_114_lpi_1_dfm_1
          | ln_land_115_lpi_1_dfm_1 | ln_land_117_lpi_1_dfm_1 | ln_land_118_lpi_1_dfm_1
          | ln_land_122_lpi_1_dfm_1 | ln_land_123_lpi_1_dfm_1 | ln_land_124_lpi_1_dfm_1
          | ln_land_125_lpi_1_dfm_1 | ln_land_126_lpi_1_dfm_1 | ln_land_132_lpi_1_dfm_1
          | ln_land_133_lpi_1_dfm_1 | ln_land_134_lpi_1_dfm_1 | ln_land_135_lpi_1_dfm_1
          | ln_land_136_lpi_1_dfm_1 | ln_land_141_lpi_1_dfm_1 | ln_land_142_lpi_1_dfm_1
          | ln_and_138_ssc_1 | ln_land_144_lpi_1_dfm_1) & (~(ln_and_140_ssc_1 | ln_land_146_lpi_1_dfm_1
          | ln_land_147_lpi_1_dfm_1 | ln_land_148_lpi_1_dfm_1 | ln_land_153_lpi_1_dfm_1
          | ln_land_154_lpi_1_dfm_1 | ln_land_155_lpi_1_dfm_1 | ln_land_156_lpi_1_dfm_1
          | ln_land_161_lpi_1_dfm_1 | ln_land_162_lpi_1_dfm_1 | ln_land_163_lpi_1_dfm_1
          | ln_land_164_lpi_1_dfm_1 | ln_land_168_lpi_1_dfm_1 | ln_land_169_lpi_1_dfm_1
          | ln_land_170_lpi_1_dfm_1 | ln_land_171_lpi_1_dfm_1 | ln_land_175_lpi_1_dfm_1
          | ln_land_176_lpi_1_dfm_1 | ln_land_177_lpi_1_dfm_1 | ln_land_181_lpi_1_dfm_1
          | ln_land_182_lpi_1_dfm_1 | ln_land_183_lpi_1_dfm_1 | ln_land_187_lpi_1_dfm_1
          | ln_land_188_lpi_1_dfm_1 | ln_land_189_lpi_1_dfm_1 | ln_land_193_lpi_1_dfm_1
          | ln_land_194_lpi_1_dfm_1 | ln_land_198_lpi_1_dfm_1 | ln_land_199_lpi_1_dfm_1
          | ln_land_200_lpi_1_dfm_1 | ln_land_203_lpi_1_dfm_1 | ln_land_204_lpi_1_dfm_1
          | ln_land_208_lpi_1_dfm_1 | ln_land_209_lpi_1_dfm_1 | ln_land_212_lpi_1_dfm_1
          | ln_land_213_lpi_1_dfm_1 | ln_land_216_lpi_1_dfm_1 | ln_land_217_lpi_1_dfm_1
          | ln_land_220_lpi_1_dfm_1 | ln_land_221_lpi_1_dfm_1 | ln_land_224_lpi_1_dfm_1
          | ln_land_227_lpi_1_dfm_1 | ln_land_228_lpi_1_dfm_1 | ln_land_230_lpi_1_dfm_1
          | ln_land_231_lpi_1_dfm_1 | ln_land_233_lpi_1_dfm_1 | ln_land_234_lpi_1_dfm_1
          | ln_land_236_lpi_1_dfm_1 | ln_land_239_lpi_1_dfm_1 | ln_land_241_lpi_1_dfm_1
          | ln_land_243_lpi_1_dfm_1))) | ln_land_149_lpi_1_dfm_1 | ln_land_150_lpi_1_dfm_1
          | ln_land_151_lpi_1_dfm_1 | ln_land_152_lpi_1_dfm_1 | ln_land_157_lpi_1_dfm_1
          | ln_land_158_lpi_1_dfm_1 | ln_land_159_lpi_1_dfm_1 | ln_land_160_lpi_1_dfm_1
          | ln_land_165_lpi_1_dfm_1 | ln_land_166_lpi_1_dfm_1 | ln_land_167_lpi_1_dfm_1
          | ln_land_172_lpi_1_dfm_1 | ln_land_173_lpi_1_dfm_1 | ln_land_174_lpi_1_dfm_1
          | ln_land_178_lpi_1_dfm_1 | ln_land_179_lpi_1_dfm_1 | ln_land_180_lpi_1_dfm_1
          | ln_land_184_lpi_1_dfm_1 | ln_land_185_lpi_1_dfm_1 | ln_land_186_lpi_1_dfm_1
          | ln_land_190_lpi_1_dfm_1 | ln_land_191_lpi_1_dfm_1 | ln_land_192_lpi_1_dfm_1
          | ln_land_195_lpi_1_dfm_1 | ln_land_196_lpi_1_dfm_1 | ln_land_197_lpi_1_dfm_1
          | ln_land_201_lpi_1_dfm_1 | ln_land_202_lpi_1_dfm_1 | ln_land_205_lpi_1_dfm_1
          | ln_land_206_lpi_1_dfm_1 | ln_land_207_lpi_1_dfm_1 | ln_land_210_lpi_1_dfm_1
          | ln_land_211_lpi_1_dfm_1 | ln_land_214_lpi_1_dfm_1 | ln_land_215_lpi_1_dfm_1
          | ln_land_218_lpi_1_dfm_1 | ln_land_219_lpi_1_dfm_1 | ln_land_222_lpi_1_dfm_1
          | ln_land_223_lpi_1_dfm_1 | ln_land_225_lpi_1_dfm_1 | ln_land_226_lpi_1_dfm_1
          | ln_land_229_lpi_1_dfm_1 | ln_land_232_lpi_1_dfm_1 | ln_land_235_lpi_1_dfm_1
          | ln_land_237_lpi_1_dfm_1 | ln_land_238_lpi_1_dfm_1 | ln_land_240_lpi_1_dfm_1
          | ln_land_242_lpi_1_dfm_1 | ln_land_244_lpi_1_dfm_1;
      ln_ln_mux1h_118_psp_1_5 <= (((((~(((~(ln_ln_ln_nor_8_cse_1 | ln_land_6_lpi_1_dfm_1
          | ln_and_2_ssc_1)) & (~(ln_and_4_ssc_1 | ln_land_8_lpi_1_dfm_1 | ln_land_12_lpi_1_dfm_1
          | ln_land_13_lpi_1_dfm_1 | ln_land_17_lpi_1_dfm_1 | ln_land_18_lpi_1_dfm_1
          | ln_land_21_lpi_1_dfm_1 | ln_land_22_lpi_1_dfm_1 | ln_land_23_lpi_1_dfm_1
          | ln_land_26_lpi_1_dfm_1 | ln_land_27_lpi_1_dfm_1 | ln_land_30_lpi_1_dfm_1
          | ln_land_31_lpi_1_dfm_1 | ln_land_35_lpi_1_dfm_1 | ln_land_36_lpi_1_dfm_1
          | ln_land_39_lpi_1_dfm_1 | ln_land_40_lpi_1_dfm_1 | ln_land_43_lpi_1_dfm_1
          | ln_land_44_lpi_1_dfm_1 | ln_land_47_lpi_1_dfm_1 | ln_land_48_lpi_1_dfm_1)))
          | ln_land_9_lpi_1_dfm_1 | ln_land_10_lpi_1_dfm_1 | ln_land_11_lpi_1_dfm_1
          | ln_land_14_lpi_1_dfm_1 | ln_land_15_lpi_1_dfm_1 | ln_land_16_lpi_1_dfm_1
          | ln_land_19_lpi_1_dfm_1 | ln_land_20_lpi_1_dfm_1 | ln_land_24_lpi_1_dfm_1
          | ln_land_25_lpi_1_dfm_1 | ln_land_28_lpi_1_dfm_1 | ln_land_29_lpi_1_dfm_1
          | ln_land_32_lpi_1_dfm_1 | ln_land_33_lpi_1_dfm_1 | ln_land_34_lpi_1_dfm_1
          | ln_land_37_lpi_1_dfm_1 | ln_land_38_lpi_1_dfm_1 | ln_land_41_lpi_1_dfm_1
          | ln_land_42_lpi_1_dfm_1 | ln_land_45_lpi_1_dfm_1 | ln_land_46_lpi_1_dfm_1
          | ln_land_49_lpi_1_dfm_1 | ln_if_50_ln_if_50_and_seb_1 | ln_land_52_lpi_1_dfm_1))
          | ln_land_51_lpi_1_dfm_1) & (~(ln_and_48_ssc_1 | ln_land_56_lpi_1_dfm_1
          | ln_land_57_lpi_1_dfm_1 | ln_land_60_lpi_1_dfm_1 | ln_land_63_lpi_1_dfm_1
          | ln_land_64_lpi_1_dfm_1 | ln_land_66_lpi_1_dfm_1 | ln_land_67_lpi_1_dfm_1
          | ln_land_69_lpi_1_dfm_1 | ln_land_70_lpi_1_dfm_1 | ln_land_73_lpi_1_dfm_1
          | ln_land_76_lpi_1_dfm_1 | ln_land_79_lpi_1_dfm_1 | ln_land_81_lpi_1_dfm_1
          | ln_land_82_lpi_1_dfm_1 | ln_land_84_lpi_1_dfm_1 | ln_land_87_lpi_1_dfm_1
          | ln_land_89_lpi_1_dfm_1 | ln_land_90_lpi_1_dfm_1 | ln_land_92_lpi_1_dfm_1
          | ln_land_94_lpi_1_dfm_1 | ln_land_97_lpi_1_dfm_1 | ln_land_99_lpi_1_dfm_1
          | ln_land_101_lpi_1_dfm_1 | ln_land_103_lpi_1_dfm_1 | ln_land_105_lpi_1_dfm_1
          | ln_land_107_lpi_1_dfm_1 | ln_land_109_lpi_1_dfm_1 | ln_land_111_lpi_1_dfm_1
          | ln_land_113_lpi_1_dfm_1 | ln_land_115_lpi_1_dfm_1 | ln_land_116_lpi_1_dfm_1
          | ln_land_118_lpi_1_dfm_1 | ln_land_120_lpi_1_dfm_1 | ln_land_121_lpi_1_dfm_1
          | ln_land_125_lpi_1_dfm_1 | ln_land_126_lpi_1_dfm_1 | ln_land_130_lpi_1_dfm_1
          | ln_land_131_lpi_1_dfm_1 | ln_land_134_lpi_1_dfm_1 | ln_land_135_lpi_1_dfm_1
          | ln_land_136_lpi_1_dfm_1 | ln_land_139_lpi_1_dfm_1 | ln_land_140_lpi_1_dfm_1)))
          | ln_land_54_lpi_1_dfm_1 | ln_land_55_lpi_1_dfm_1 | ln_land_58_lpi_1_dfm_1
          | ln_land_59_lpi_1_dfm_1 | ln_land_61_lpi_1_dfm_1 | ln_land_62_lpi_1_dfm_1
          | ln_land_65_lpi_1_dfm_1 | ln_land_68_lpi_1_dfm_1 | ln_land_71_lpi_1_dfm_1
          | ln_land_72_lpi_1_dfm_1 | ln_land_74_lpi_1_dfm_1 | ln_land_75_lpi_1_dfm_1
          | ln_land_77_lpi_1_dfm_1 | ln_land_78_lpi_1_dfm_1 | ln_land_80_lpi_1_dfm_1
          | ln_land_83_lpi_1_dfm_1 | ln_land_85_lpi_1_dfm_1 | ln_land_86_lpi_1_dfm_1
          | ln_land_88_lpi_1_dfm_1 | ln_land_91_lpi_1_dfm_1 | ln_land_93_lpi_1_dfm_1
          | ln_land_95_lpi_1_dfm_1 | ln_land_96_lpi_1_dfm_1 | ln_land_98_lpi_1_dfm_1
          | ln_land_100_lpi_1_dfm_1 | ln_land_102_lpi_1_dfm_1 | ln_land_104_lpi_1_dfm_1
          | ln_land_106_lpi_1_dfm_1 | ln_land_108_lpi_1_dfm_1 | ln_land_110_lpi_1_dfm_1
          | ln_land_112_lpi_1_dfm_1 | ln_land_114_lpi_1_dfm_1 | ln_land_117_lpi_1_dfm_1
          | ln_land_119_lpi_1_dfm_1 | ln_land_122_lpi_1_dfm_1 | ln_land_123_lpi_1_dfm_1
          | ln_land_124_lpi_1_dfm_1 | ln_land_127_lpi_1_dfm_1 | ln_land_128_lpi_1_dfm_1
          | ln_land_129_lpi_1_dfm_1 | ln_land_132_lpi_1_dfm_1 | ln_land_133_lpi_1_dfm_1
          | ln_land_137_lpi_1_dfm_1 | ln_land_138_lpi_1_dfm_1 | ln_land_141_lpi_1_dfm_1
          | ln_land_142_lpi_1_dfm_1) & ln_nor_3_cse_1 & (~(ln_land_147_lpi_1_dfm_1
          | ln_land_148_lpi_1_dfm_1 | ln_land_151_lpi_1_dfm_1 | ln_land_152_lpi_1_dfm_1
          | ln_land_155_lpi_1_dfm_1 | ln_land_156_lpi_1_dfm_1 | ln_land_159_lpi_1_dfm_1
          | ln_land_160_lpi_1_dfm_1 | ln_land_163_lpi_1_dfm_1 | ln_land_164_lpi_1_dfm_1
          | ln_land_166_lpi_1_dfm_1 | ln_land_167_lpi_1_dfm_1 | ln_land_170_lpi_1_dfm_1
          | ln_land_171_lpi_1_dfm_1 | ln_land_173_lpi_1_dfm_1 | ln_land_174_lpi_1_dfm_1
          | ln_land_177_lpi_1_dfm_1 | ln_land_180_lpi_1_dfm_1 | ln_land_183_lpi_1_dfm_1
          | ln_land_186_lpi_1_dfm_1 | ln_land_189_lpi_1_dfm_1 | ln_land_191_lpi_1_dfm_1
          | ln_land_192_lpi_1_dfm_1 | ln_land_194_lpi_1_dfm_1 | ln_land_197_lpi_1_dfm_1
          | ln_land_199_lpi_1_dfm_1 | ln_land_200_lpi_1_dfm_1 | ln_land_202_lpi_1_dfm_1
          | ln_land_204_lpi_1_dfm_1 | ln_land_206_lpi_1_dfm_1 | ln_land_207_lpi_1_dfm_1
          | ln_land_209_lpi_1_dfm_1 | ln_land_211_lpi_1_dfm_1 | ln_land_213_lpi_1_dfm_1
          | ln_land_215_lpi_1_dfm_1 | ln_land_217_lpi_1_dfm_1 | ln_land_219_lpi_1_dfm_1
          | ln_land_221_lpi_1_dfm_1 | ln_land_223_lpi_1_dfm_1 | ln_land_224_lpi_1_dfm_1
          | ln_land_226_lpi_1_dfm_1 | ln_land_228_lpi_1_dfm_1 | ln_land_229_lpi_1_dfm_1
          | ln_land_231_lpi_1_dfm_1 | ln_land_232_lpi_1_dfm_1 | ln_land_234_lpi_1_dfm_1
          | ln_land_235_lpi_1_dfm_1 | ln_land_238_lpi_1_dfm_1 | ln_land_239_lpi_1_dfm_1
          | ln_land_240_lpi_1_dfm_1))) | ln_and_140_ssc_1 | ln_land_146_lpi_1_dfm_1
          | ln_land_149_lpi_1_dfm_1 | ln_land_150_lpi_1_dfm_1 | ln_land_153_lpi_1_dfm_1
          | ln_land_154_lpi_1_dfm_1 | ln_land_157_lpi_1_dfm_1 | ln_land_158_lpi_1_dfm_1
          | ln_land_161_lpi_1_dfm_1 | ln_land_162_lpi_1_dfm_1 | ln_land_165_lpi_1_dfm_1
          | ln_land_168_lpi_1_dfm_1 | ln_land_169_lpi_1_dfm_1 | ln_land_172_lpi_1_dfm_1
          | ln_land_175_lpi_1_dfm_1 | ln_land_176_lpi_1_dfm_1 | ln_land_178_lpi_1_dfm_1
          | ln_land_179_lpi_1_dfm_1 | ln_land_181_lpi_1_dfm_1 | ln_land_182_lpi_1_dfm_1
          | ln_land_184_lpi_1_dfm_1 | ln_land_185_lpi_1_dfm_1 | ln_land_187_lpi_1_dfm_1
          | ln_land_188_lpi_1_dfm_1 | ln_land_190_lpi_1_dfm_1 | ln_land_193_lpi_1_dfm_1
          | ln_land_195_lpi_1_dfm_1 | ln_land_196_lpi_1_dfm_1 | ln_land_198_lpi_1_dfm_1
          | ln_land_201_lpi_1_dfm_1 | ln_land_203_lpi_1_dfm_1 | ln_land_205_lpi_1_dfm_1
          | ln_land_208_lpi_1_dfm_1 | ln_land_210_lpi_1_dfm_1 | ln_land_212_lpi_1_dfm_1
          | ln_land_214_lpi_1_dfm_1 | ln_land_216_lpi_1_dfm_1 | ln_land_218_lpi_1_dfm_1
          | ln_land_220_lpi_1_dfm_1 | ln_land_222_lpi_1_dfm_1 | ln_land_225_lpi_1_dfm_1
          | ln_land_227_lpi_1_dfm_1 | ln_land_230_lpi_1_dfm_1 | ln_land_233_lpi_1_dfm_1
          | ln_land_236_lpi_1_dfm_1 | ln_land_237_lpi_1_dfm_1 | ln_land_241_lpi_1_dfm_1
          | ln_land_242_lpi_1_dfm_1 | ln_land_243_lpi_1_dfm_1 | ln_land_244_lpi_1_dfm_1;
      ln_ln_mux1h_118_psp_1_4 <= (((~((~((~((~((((~(((~((~((~(ln_ret_13_0_lpi_1_dfm_258
          | ln_land_3_lpi_1_dfm_1)) | ln_land_4_lpi_1_dfm_1 | ln_land_6_lpi_1_dfm_1))
          | ln_and_2_ssc_1)) & (~(ln_and_4_ssc_1 | ln_land_9_lpi_1_dfm_1 | ln_land_12_lpi_1_dfm_1
          | ln_land_14_lpi_1_dfm_1 | ln_land_17_lpi_1_dfm_1 | ln_land_19_lpi_1_dfm_1
          | ln_land_21_lpi_1_dfm_1 | ln_land_24_lpi_1_dfm_1 | ln_land_26_lpi_1_dfm_1
          | ln_land_28_lpi_1_dfm_1 | ln_land_30_lpi_1_dfm_1 | ln_land_32_lpi_1_dfm_1
          | ln_land_33_lpi_1_dfm_1 | ln_land_35_lpi_1_dfm_1 | ln_land_37_lpi_1_dfm_1
          | ln_land_39_lpi_1_dfm_1 | ln_land_41_lpi_1_dfm_1 | ln_land_43_lpi_1_dfm_1
          | ln_land_45_lpi_1_dfm_1 | ln_land_47_lpi_1_dfm_1 | ln_land_49_lpi_1_dfm_1)))
          | ln_land_8_lpi_1_dfm_1 | ln_land_10_lpi_1_dfm_1 | ln_land_11_lpi_1_dfm_1
          | ln_land_13_lpi_1_dfm_1 | ln_land_15_lpi_1_dfm_1 | ln_land_16_lpi_1_dfm_1
          | ln_land_18_lpi_1_dfm_1 | ln_land_20_lpi_1_dfm_1 | ln_land_22_lpi_1_dfm_1
          | ln_land_23_lpi_1_dfm_1 | ln_land_25_lpi_1_dfm_1 | ln_land_27_lpi_1_dfm_1
          | ln_land_29_lpi_1_dfm_1 | ln_land_31_lpi_1_dfm_1 | ln_land_34_lpi_1_dfm_1
          | ln_land_36_lpi_1_dfm_1 | ln_land_38_lpi_1_dfm_1 | ln_land_40_lpi_1_dfm_1
          | ln_land_42_lpi_1_dfm_1 | ln_land_44_lpi_1_dfm_1 | ln_land_46_lpi_1_dfm_1
          | ln_land_48_lpi_1_dfm_1 | ln_if_50_ln_if_50_and_seb_1 | ln_land_51_lpi_1_dfm_1))
          | ln_land_52_lpi_1_dfm_1) & (~(ln_and_48_ssc_1 | ln_land_55_lpi_1_dfm_1
          | ln_land_57_lpi_1_dfm_1 | ln_land_59_lpi_1_dfm_1 | ln_land_60_lpi_1_dfm_1
          | ln_land_62_lpi_1_dfm_1 | ln_land_64_lpi_1_dfm_1 | ln_land_65_lpi_1_dfm_1
          | ln_land_67_lpi_1_dfm_1 | ln_land_70_lpi_1_dfm_1 | ln_land_72_lpi_1_dfm_1
          | ln_land_73_lpi_1_dfm_1 | ln_land_75_lpi_1_dfm_1 | ln_land_76_lpi_1_dfm_1
          | ln_land_78_lpi_1_dfm_1 | ln_land_79_lpi_1_dfm_1 | ln_land_82_lpi_1_dfm_1
          | ln_land_83_lpi_1_dfm_1 | ln_land_86_lpi_1_dfm_1 | ln_land_87_lpi_1_dfm_1
          | ln_land_90_lpi_1_dfm_1 | ln_land_91_lpi_1_dfm_1 | ln_land_92_lpi_1_dfm_1
          | ln_land_96_lpi_1_dfm_1 | ln_land_97_lpi_1_dfm_1 | ln_land_98_lpi_1_dfm_1
          | ln_land_99_lpi_1_dfm_1 | ln_land_100_lpi_1_dfm_1 | ln_land_112_lpi_1_dfm_1
          | ln_land_113_lpi_1_dfm_1 | ln_land_114_lpi_1_dfm_1 | ln_land_115_lpi_1_dfm_1
          | ln_land_118_lpi_1_dfm_1 | ln_land_119_lpi_1_dfm_1 | ln_land_121_lpi_1_dfm_1
          | ln_land_124_lpi_1_dfm_1 | ln_land_126_lpi_1_dfm_1 | ln_land_128_lpi_1_dfm_1
          | ln_land_129_lpi_1_dfm_1 | ln_land_131_lpi_1_dfm_1 | ln_land_133_lpi_1_dfm_1
          | ln_land_135_lpi_1_dfm_1 | ln_land_136_lpi_1_dfm_1 | ln_land_138_lpi_1_dfm_1
          | ln_land_140_lpi_1_dfm_1))) | ln_land_54_lpi_1_dfm_1 | ln_land_56_lpi_1_dfm_1
          | ln_land_58_lpi_1_dfm_1 | ln_land_61_lpi_1_dfm_1 | ln_land_63_lpi_1_dfm_1
          | ln_land_66_lpi_1_dfm_1 | ln_land_68_lpi_1_dfm_1 | ln_land_69_lpi_1_dfm_1
          | ln_land_71_lpi_1_dfm_1 | ln_land_74_lpi_1_dfm_1 | ln_land_77_lpi_1_dfm_1
          | ln_land_80_lpi_1_dfm_1 | ln_land_81_lpi_1_dfm_1 | ln_land_84_lpi_1_dfm_1
          | ln_land_85_lpi_1_dfm_1 | ln_land_88_lpi_1_dfm_1 | ln_land_89_lpi_1_dfm_1
          | ln_land_93_lpi_1_dfm_1 | ln_land_94_lpi_1_dfm_1 | ln_land_95_lpi_1_dfm_1
          | ln_land_101_lpi_1_dfm_1 | ln_land_102_lpi_1_dfm_1 | ln_land_103_lpi_1_dfm_1
          | ln_land_104_lpi_1_dfm_1 | ln_land_105_lpi_1_dfm_1 | ln_land_106_lpi_1_dfm_1
          | ln_land_107_lpi_1_dfm_1 | ln_land_108_lpi_1_dfm_1 | ln_land_109_lpi_1_dfm_1
          | ln_land_110_lpi_1_dfm_1 | ln_land_111_lpi_1_dfm_1 | ln_land_116_lpi_1_dfm_1
          | ln_land_117_lpi_1_dfm_1 | ln_land_120_lpi_1_dfm_1 | ln_land_122_lpi_1_dfm_1
          | ln_land_123_lpi_1_dfm_1 | ln_land_125_lpi_1_dfm_1 | ln_land_127_lpi_1_dfm_1
          | ln_land_130_lpi_1_dfm_1 | ln_land_132_lpi_1_dfm_1 | ln_land_134_lpi_1_dfm_1
          | ln_land_137_lpi_1_dfm_1 | ln_land_139_lpi_1_dfm_1)) | ln_land_142_lpi_1_dfm_1))
          | ln_land_141_lpi_1_dfm_1)) | ln_land_144_lpi_1_dfm_1)) | ln_and_138_ssc_1)
          & (~(ln_land_146_lpi_1_dfm_1 | ln_land_148_lpi_1_dfm_1 | ln_land_150_lpi_1_dfm_1
          | ln_land_152_lpi_1_dfm_1 | ln_land_154_lpi_1_dfm_1 | ln_land_156_lpi_1_dfm_1
          | ln_land_158_lpi_1_dfm_1 | ln_land_160_lpi_1_dfm_1 | ln_land_162_lpi_1_dfm_1
          | ln_land_164_lpi_1_dfm_1 | ln_land_167_lpi_1_dfm_1 | ln_land_169_lpi_1_dfm_1
          | ln_land_171_lpi_1_dfm_1 | ln_land_172_lpi_1_dfm_1 | ln_land_174_lpi_1_dfm_1
          | ln_land_176_lpi_1_dfm_1 | ln_land_177_lpi_1_dfm_1 | ln_land_179_lpi_1_dfm_1
          | ln_land_180_lpi_1_dfm_1 | ln_land_182_lpi_1_dfm_1 | ln_land_185_lpi_1_dfm_1
          | ln_land_186_lpi_1_dfm_1 | ln_land_188_lpi_1_dfm_1 | ln_land_189_lpi_1_dfm_1
          | ln_land_192_lpi_1_dfm_1 | ln_land_193_lpi_1_dfm_1 | ln_land_196_lpi_1_dfm_1
          | ln_land_197_lpi_1_dfm_1 | ln_land_200_lpi_1_dfm_1 | ln_land_201_lpi_1_dfm_1
          | ln_land_202_lpi_1_dfm_1 | ln_land_207_lpi_1_dfm_1 | ln_land_208_lpi_1_dfm_1
          | ln_land_209_lpi_1_dfm_1 | ln_land_210_lpi_1_dfm_1 | ln_land_211_lpi_1_dfm_1
          | ln_land_212_lpi_1_dfm_1 | ln_land_218_lpi_1_dfm_1 | ln_land_219_lpi_1_dfm_1
          | ln_land_220_lpi_1_dfm_1 | ln_land_221_lpi_1_dfm_1 | ln_land_222_lpi_1_dfm_1
          | ln_land_223_lpi_1_dfm_1 | ln_land_226_lpi_1_dfm_1 | ln_land_227_lpi_1_dfm_1
          | ln_land_228_lpi_1_dfm_1 | ln_land_230_lpi_1_dfm_1 | ln_land_231_lpi_1_dfm_1
          | ln_land_233_lpi_1_dfm_1 | ln_land_234_lpi_1_dfm_1 | ln_land_236_lpi_1_dfm_1
          | ln_land_238_lpi_1_dfm_1 | ln_land_239_lpi_1_dfm_1 | ln_land_241_lpi_1_dfm_1
          | ln_land_242_lpi_1_dfm_1))) | ln_and_140_ssc_1 | ln_land_147_lpi_1_dfm_1
          | ln_land_149_lpi_1_dfm_1 | ln_land_151_lpi_1_dfm_1 | ln_land_153_lpi_1_dfm_1
          | ln_land_155_lpi_1_dfm_1 | ln_land_157_lpi_1_dfm_1 | ln_land_159_lpi_1_dfm_1
          | ln_land_161_lpi_1_dfm_1 | ln_land_163_lpi_1_dfm_1 | ln_land_165_lpi_1_dfm_1
          | ln_land_166_lpi_1_dfm_1 | ln_land_168_lpi_1_dfm_1 | ln_land_170_lpi_1_dfm_1
          | ln_land_173_lpi_1_dfm_1 | ln_land_175_lpi_1_dfm_1 | ln_land_178_lpi_1_dfm_1
          | ln_land_181_lpi_1_dfm_1 | ln_land_183_lpi_1_dfm_1 | ln_land_184_lpi_1_dfm_1
          | ln_land_187_lpi_1_dfm_1 | ln_land_190_lpi_1_dfm_1 | ln_land_191_lpi_1_dfm_1
          | ln_land_194_lpi_1_dfm_1 | ln_land_195_lpi_1_dfm_1 | ln_land_198_lpi_1_dfm_1
          | ln_land_199_lpi_1_dfm_1 | ln_land_203_lpi_1_dfm_1 | ln_land_204_lpi_1_dfm_1
          | ln_land_205_lpi_1_dfm_1 | ln_land_206_lpi_1_dfm_1 | ln_land_213_lpi_1_dfm_1
          | ln_land_214_lpi_1_dfm_1 | ln_land_215_lpi_1_dfm_1 | ln_land_216_lpi_1_dfm_1
          | ln_land_217_lpi_1_dfm_1 | ln_land_224_lpi_1_dfm_1 | ln_land_225_lpi_1_dfm_1
          | ln_land_229_lpi_1_dfm_1 | ln_land_232_lpi_1_dfm_1 | ln_land_235_lpi_1_dfm_1
          | ln_land_237_lpi_1_dfm_1 | ln_land_240_lpi_1_dfm_1 | ln_land_243_lpi_1_dfm_1
          | ln_land_244_lpi_1_dfm_1;
      ln_ln_mux1h_118_psp_1_3 <= (((~((~((((~(((~((~(ln_ret_13_0_lpi_1_dfm_258 |
          ln_land_3_lpi_1_dfm_1 | ln_land_4_lpi_1_dfm_1 | ln_land_6_lpi_1_dfm_1))
          | ln_and_2_ssc_1)) & (~(ln_land_9_lpi_1_dfm_1 | ln_land_10_lpi_1_dfm_1
          | ln_land_14_lpi_1_dfm_1 | ln_land_15_lpi_1_dfm_1 | ln_land_20_lpi_1_dfm_1
          | ln_land_21_lpi_1_dfm_1 | ln_land_22_lpi_1_dfm_1 | ln_land_27_lpi_1_dfm_1
          | ln_land_28_lpi_1_dfm_1 | ln_land_29_lpi_1_dfm_1 | ln_land_30_lpi_1_dfm_1
          | ln_land_31_lpi_1_dfm_1 | ln_land_32_lpi_1_dfm_1))) | ln_and_4_ssc_1 |
          ln_land_8_lpi_1_dfm_1 | ln_land_11_lpi_1_dfm_1 | ln_land_12_lpi_1_dfm_1
          | ln_land_13_lpi_1_dfm_1 | ln_land_16_lpi_1_dfm_1 | ln_land_17_lpi_1_dfm_1
          | ln_land_18_lpi_1_dfm_1 | ln_land_19_lpi_1_dfm_1 | ln_land_23_lpi_1_dfm_1
          | ln_land_24_lpi_1_dfm_1 | ln_land_25_lpi_1_dfm_1 | ln_land_26_lpi_1_dfm_1
          | ln_land_33_lpi_1_dfm_1 | ln_land_34_lpi_1_dfm_1 | ln_land_35_lpi_1_dfm_1
          | ln_land_36_lpi_1_dfm_1 | ln_land_37_lpi_1_dfm_1 | ln_land_38_lpi_1_dfm_1
          | ln_land_39_lpi_1_dfm_1 | ln_land_40_lpi_1_dfm_1 | ln_land_41_lpi_1_dfm_1
          | ln_land_42_lpi_1_dfm_1 | ln_land_43_lpi_1_dfm_1 | ln_land_44_lpi_1_dfm_1
          | ln_land_45_lpi_1_dfm_1 | ln_land_46_lpi_1_dfm_1 | ln_land_47_lpi_1_dfm_1
          | ln_land_48_lpi_1_dfm_1 | ln_land_49_lpi_1_dfm_1 | ln_if_50_ln_if_50_and_seb_1))
          | ln_land_51_lpi_1_dfm_1 | ln_land_52_lpi_1_dfm_1) & (~(ln_land_56_lpi_1_dfm_1
          | ln_land_57_lpi_1_dfm_1 | ln_land_58_lpi_1_dfm_1 | ln_land_59_lpi_1_dfm_1
          | ln_land_63_lpi_1_dfm_1 | ln_land_64_lpi_1_dfm_1 | ln_land_67_lpi_1_dfm_1
          | ln_land_68_lpi_1_dfm_1 | ln_land_71_lpi_1_dfm_1 | ln_land_72_lpi_1_dfm_1
          | ln_land_74_lpi_1_dfm_1 | ln_land_75_lpi_1_dfm_1 | ln_land_77_lpi_1_dfm_1
          | ln_land_78_lpi_1_dfm_1 | ln_land_80_lpi_1_dfm_1 | ln_land_82_lpi_1_dfm_1
          | ln_land_84_lpi_1_dfm_1 | ln_land_86_lpi_1_dfm_1 | ln_land_88_lpi_1_dfm_1
          | ln_land_90_lpi_1_dfm_1 | ln_land_91_lpi_1_dfm_1 | ln_land_93_lpi_1_dfm_1
          | ln_land_96_lpi_1_dfm_1 | ln_land_97_lpi_1_dfm_1 | ln_land_101_lpi_1_dfm_1
          | ln_land_102_lpi_1_dfm_1 | ln_land_103_lpi_1_dfm_1 | ln_land_104_lpi_1_dfm_1
          | ln_land_105_lpi_1_dfm_1 | ln_land_107_lpi_1_dfm_1 | ln_land_108_lpi_1_dfm_1
          | ln_land_109_lpi_1_dfm_1 | ln_land_110_lpi_1_dfm_1 | ln_land_111_lpi_1_dfm_1
          | ln_land_114_lpi_1_dfm_1 | ln_land_115_lpi_1_dfm_1 | ln_land_117_lpi_1_dfm_1
          | ln_land_119_lpi_1_dfm_1 | ln_land_123_lpi_1_dfm_1 | ln_land_124_lpi_1_dfm_1
          | ln_land_129_lpi_1_dfm_1 | ln_land_130_lpi_1_dfm_1 | ln_land_131_lpi_1_dfm_1
          | ln_land_136_lpi_1_dfm_1 | ln_land_137_lpi_1_dfm_1 | ln_land_138_lpi_1_dfm_1
          | ln_land_139_lpi_1_dfm_1 | ln_land_140_lpi_1_dfm_1))) | ln_and_48_ssc_1
          | ln_land_54_lpi_1_dfm_1 | ln_land_55_lpi_1_dfm_1 | ln_land_60_lpi_1_dfm_1
          | ln_land_61_lpi_1_dfm_1 | ln_land_62_lpi_1_dfm_1 | ln_land_65_lpi_1_dfm_1
          | ln_land_66_lpi_1_dfm_1 | ln_land_69_lpi_1_dfm_1 | ln_land_70_lpi_1_dfm_1
          | ln_land_73_lpi_1_dfm_1 | ln_land_76_lpi_1_dfm_1 | ln_land_79_lpi_1_dfm_1
          | ln_land_81_lpi_1_dfm_1 | ln_land_83_lpi_1_dfm_1 | ln_land_85_lpi_1_dfm_1
          | ln_land_87_lpi_1_dfm_1 | ln_land_89_lpi_1_dfm_1 | ln_land_92_lpi_1_dfm_1
          | ln_land_94_lpi_1_dfm_1 | ln_land_95_lpi_1_dfm_1 | ln_land_98_lpi_1_dfm_1
          | ln_land_99_lpi_1_dfm_1 | ln_land_100_lpi_1_dfm_1 | ln_land_106_lpi_1_dfm_1
          | ln_land_112_lpi_1_dfm_1 | ln_land_113_lpi_1_dfm_1 | ln_land_116_lpi_1_dfm_1
          | ln_land_118_lpi_1_dfm_1 | ln_land_120_lpi_1_dfm_1 | ln_land_121_lpi_1_dfm_1
          | ln_land_122_lpi_1_dfm_1 | ln_land_125_lpi_1_dfm_1 | ln_land_126_lpi_1_dfm_1
          | ln_land_127_lpi_1_dfm_1 | ln_land_128_lpi_1_dfm_1 | ln_land_132_lpi_1_dfm_1
          | ln_land_133_lpi_1_dfm_1 | ln_land_134_lpi_1_dfm_1 | ln_land_135_lpi_1_dfm_1))
          | ln_land_141_lpi_1_dfm_1)) | ln_land_142_lpi_1_dfm_1 | ln_and_138_ssc_1
          | ln_land_144_lpi_1_dfm_1) & (~(ln_land_160_lpi_1_dfm_1 | ln_land_161_lpi_1_dfm_1
          | ln_land_162_lpi_1_dfm_1 | ln_land_163_lpi_1_dfm_1 | ln_land_164_lpi_1_dfm_1
          | ln_land_165_lpi_1_dfm_1 | ln_land_169_lpi_1_dfm_1 | ln_land_170_lpi_1_dfm_1
          | ln_land_171_lpi_1_dfm_1 | ln_land_174_lpi_1_dfm_1 | ln_land_175_lpi_1_dfm_1
          | ln_land_176_lpi_1_dfm_1 | ln_land_179_lpi_1_dfm_1 | ln_land_182_lpi_1_dfm_1
          | ln_land_183_lpi_1_dfm_1 | ln_land_185_lpi_1_dfm_1 | ln_land_188_lpi_1_dfm_1
          | ln_land_190_lpi_1_dfm_1 | ln_land_192_lpi_1_dfm_1 | ln_land_194_lpi_1_dfm_1
          | ln_land_196_lpi_1_dfm_1 | ln_land_198_lpi_1_dfm_1 | ln_land_200_lpi_1_dfm_1
          | ln_land_201_lpi_1_dfm_1 | ln_land_203_lpi_1_dfm_1 | ln_land_204_lpi_1_dfm_1
          | ln_land_207_lpi_1_dfm_1 | ln_land_208_lpi_1_dfm_1 | ln_land_213_lpi_1_dfm_1
          | ln_land_214_lpi_1_dfm_1 | ln_land_215_lpi_1_dfm_1 | ln_land_216_lpi_1_dfm_1
          | ln_land_217_lpi_1_dfm_1 | ln_land_222_lpi_1_dfm_1 | ln_land_223_lpi_1_dfm_1
          | ln_land_225_lpi_1_dfm_1 | ln_land_228_lpi_1_dfm_1 | ln_land_231_lpi_1_dfm_1
          | ln_land_234_lpi_1_dfm_1 | ln_land_235_lpi_1_dfm_1 | ln_land_236_lpi_1_dfm_1
          | ln_land_237_lpi_1_dfm_1 | ln_land_238_lpi_1_dfm_1 | ln_land_241_lpi_1_dfm_1
          | ln_land_243_lpi_1_dfm_1))) | ln_and_140_ssc_1 | ln_land_146_lpi_1_dfm_1
          | ln_land_147_lpi_1_dfm_1 | ln_land_148_lpi_1_dfm_1 | ln_land_149_lpi_1_dfm_1
          | ln_land_150_lpi_1_dfm_1 | ln_land_151_lpi_1_dfm_1 | ln_land_152_lpi_1_dfm_1
          | ln_land_153_lpi_1_dfm_1 | ln_land_154_lpi_1_dfm_1 | ln_land_155_lpi_1_dfm_1
          | ln_land_156_lpi_1_dfm_1 | ln_land_157_lpi_1_dfm_1 | ln_land_158_lpi_1_dfm_1
          | ln_land_159_lpi_1_dfm_1 | ln_land_166_lpi_1_dfm_1 | ln_land_167_lpi_1_dfm_1
          | ln_land_168_lpi_1_dfm_1 | ln_land_172_lpi_1_dfm_1 | ln_land_173_lpi_1_dfm_1
          | ln_land_177_lpi_1_dfm_1 | ln_land_178_lpi_1_dfm_1 | ln_land_180_lpi_1_dfm_1
          | ln_land_181_lpi_1_dfm_1 | ln_land_184_lpi_1_dfm_1 | ln_land_186_lpi_1_dfm_1
          | ln_land_187_lpi_1_dfm_1 | ln_land_189_lpi_1_dfm_1 | ln_land_191_lpi_1_dfm_1
          | ln_land_193_lpi_1_dfm_1 | ln_land_195_lpi_1_dfm_1 | ln_land_197_lpi_1_dfm_1
          | ln_land_199_lpi_1_dfm_1 | ln_land_202_lpi_1_dfm_1 | ln_land_205_lpi_1_dfm_1
          | ln_land_206_lpi_1_dfm_1 | ln_land_209_lpi_1_dfm_1 | ln_land_210_lpi_1_dfm_1
          | ln_land_211_lpi_1_dfm_1 | ln_land_212_lpi_1_dfm_1 | ln_land_218_lpi_1_dfm_1
          | ln_land_219_lpi_1_dfm_1 | ln_land_220_lpi_1_dfm_1 | ln_land_221_lpi_1_dfm_1
          | ln_land_224_lpi_1_dfm_1 | ln_land_226_lpi_1_dfm_1 | ln_land_227_lpi_1_dfm_1
          | ln_land_229_lpi_1_dfm_1 | ln_land_230_lpi_1_dfm_1 | ln_land_232_lpi_1_dfm_1
          | ln_land_233_lpi_1_dfm_1 | ln_land_239_lpi_1_dfm_1 | ln_land_240_lpi_1_dfm_1
          | ln_land_242_lpi_1_dfm_1 | ln_land_244_lpi_1_dfm_1;
      ln_ln_mux1h_118_psp_1_2 <= (((~((~((((~(((~(ln_nor_5_cse_1 | ln_and_2_ssc_1
          | ln_land_6_lpi_1_dfm_1)) & (~(ln_and_4_ssc_1 | ln_land_8_lpi_1_dfm_1 |
          ln_land_10_lpi_1_dfm_1 | ln_land_12_lpi_1_dfm_1 | ln_land_13_lpi_1_dfm_1
          | ln_land_15_lpi_1_dfm_1 | ln_land_18_lpi_1_dfm_1 | ln_land_19_lpi_1_dfm_1
          | ln_land_21_lpi_1_dfm_1 | ln_land_22_lpi_1_dfm_1 | ln_land_25_lpi_1_dfm_1
          | ln_land_26_lpi_1_dfm_1 | ln_land_30_lpi_1_dfm_1 | ln_land_31_lpi_1_dfm_1
          | ln_land_32_lpi_1_dfm_1 | ln_land_38_lpi_1_dfm_1 | ln_land_39_lpi_1_dfm_1
          | ln_land_40_lpi_1_dfm_1 | ln_land_41_lpi_1_dfm_1 | ln_land_42_lpi_1_dfm_1
          | ln_land_43_lpi_1_dfm_1 | ln_land_44_lpi_1_dfm_1 | ln_land_45_lpi_1_dfm_1
          | ln_land_46_lpi_1_dfm_1))) | ln_land_9_lpi_1_dfm_1 | ln_land_11_lpi_1_dfm_1
          | ln_land_14_lpi_1_dfm_1 | ln_land_16_lpi_1_dfm_1 | ln_land_17_lpi_1_dfm_1
          | ln_land_20_lpi_1_dfm_1 | ln_land_23_lpi_1_dfm_1 | ln_land_24_lpi_1_dfm_1
          | ln_land_27_lpi_1_dfm_1 | ln_land_28_lpi_1_dfm_1 | ln_land_29_lpi_1_dfm_1
          | ln_land_33_lpi_1_dfm_1 | ln_land_34_lpi_1_dfm_1 | ln_land_35_lpi_1_dfm_1
          | ln_land_36_lpi_1_dfm_1 | ln_land_37_lpi_1_dfm_1 | ln_land_47_lpi_1_dfm_1
          | ln_land_48_lpi_1_dfm_1 | ln_land_49_lpi_1_dfm_1 | ln_if_50_ln_if_50_and_seb_1))
          | ln_land_51_lpi_1_dfm_1 | ln_land_52_lpi_1_dfm_1) & (~(ln_land_54_lpi_1_dfm_1
          | ln_land_55_lpi_1_dfm_1 | ln_land_58_lpi_1_dfm_1 | ln_land_59_lpi_1_dfm_1
          | ln_land_61_lpi_1_dfm_1 | ln_land_62_lpi_1_dfm_1 | ln_land_64_lpi_1_dfm_1
          | ln_land_66_lpi_1_dfm_1 | ln_land_68_lpi_1_dfm_1 | ln_land_70_lpi_1_dfm_1
          | ln_land_72_lpi_1_dfm_1 | ln_land_75_lpi_1_dfm_1 | ln_land_78_lpi_1_dfm_1
          | ln_land_79_lpi_1_dfm_1 | ln_land_80_lpi_1_dfm_1 | ln_land_89_lpi_1_dfm_1
          | ln_land_90_lpi_1_dfm_1 | ln_land_93_lpi_1_dfm_1 | ln_land_94_lpi_1_dfm_1
          | ln_land_96_lpi_1_dfm_1 | ln_land_98_lpi_1_dfm_1 | ln_land_101_lpi_1_dfm_1
          | ln_land_106_lpi_1_dfm_1 | ln_land_110_lpi_1_dfm_1 | ln_land_111_lpi_1_dfm_1
          | ln_land_113_lpi_1_dfm_1 | ln_land_115_lpi_1_dfm_1 | ln_land_116_lpi_1_dfm_1
          | ln_land_120_lpi_1_dfm_1 | ln_land_123_lpi_1_dfm_1 | ln_land_125_lpi_1_dfm_1
          | ln_land_126_lpi_1_dfm_1 | ln_land_129_lpi_1_dfm_1 | ln_land_132_lpi_1_dfm_1
          | ln_land_133_lpi_1_dfm_1 | ln_land_136_lpi_1_dfm_1 | ln_land_137_lpi_1_dfm_1
          | ln_land_138_lpi_1_dfm_1))) | ln_and_48_ssc_1 | ln_land_56_lpi_1_dfm_1
          | ln_land_57_lpi_1_dfm_1 | ln_land_60_lpi_1_dfm_1 | ln_land_63_lpi_1_dfm_1
          | ln_land_65_lpi_1_dfm_1 | ln_land_67_lpi_1_dfm_1 | ln_land_69_lpi_1_dfm_1
          | ln_land_71_lpi_1_dfm_1 | ln_land_73_lpi_1_dfm_1 | ln_land_74_lpi_1_dfm_1
          | ln_land_76_lpi_1_dfm_1 | ln_land_77_lpi_1_dfm_1 | ln_land_81_lpi_1_dfm_1
          | ln_land_82_lpi_1_dfm_1 | ln_land_83_lpi_1_dfm_1 | ln_land_84_lpi_1_dfm_1
          | ln_land_85_lpi_1_dfm_1 | ln_land_86_lpi_1_dfm_1 | ln_land_87_lpi_1_dfm_1
          | ln_land_88_lpi_1_dfm_1 | ln_land_91_lpi_1_dfm_1 | ln_land_92_lpi_1_dfm_1
          | ln_land_95_lpi_1_dfm_1 | ln_land_97_lpi_1_dfm_1 | ln_land_99_lpi_1_dfm_1
          | ln_land_100_lpi_1_dfm_1 | ln_land_102_lpi_1_dfm_1 | ln_land_103_lpi_1_dfm_1
          | ln_land_104_lpi_1_dfm_1 | ln_land_105_lpi_1_dfm_1 | ln_land_107_lpi_1_dfm_1
          | ln_land_108_lpi_1_dfm_1 | ln_land_109_lpi_1_dfm_1 | ln_land_112_lpi_1_dfm_1
          | ln_land_114_lpi_1_dfm_1 | ln_land_117_lpi_1_dfm_1 | ln_land_118_lpi_1_dfm_1
          | ln_land_119_lpi_1_dfm_1 | ln_land_121_lpi_1_dfm_1 | ln_land_122_lpi_1_dfm_1
          | ln_land_124_lpi_1_dfm_1 | ln_land_127_lpi_1_dfm_1 | ln_land_128_lpi_1_dfm_1
          | ln_land_130_lpi_1_dfm_1 | ln_land_131_lpi_1_dfm_1 | ln_land_134_lpi_1_dfm_1
          | ln_land_135_lpi_1_dfm_1 | ln_land_139_lpi_1_dfm_1 | ln_land_140_lpi_1_dfm_1))
          | ln_land_142_lpi_1_dfm_1)) | ln_land_141_lpi_1_dfm_1) & ln_nor_3_cse_1
          & (~(ln_and_140_ssc_1 | ln_land_146_lpi_1_dfm_1 | ln_land_156_lpi_1_dfm_1
          | ln_land_157_lpi_1_dfm_1 | ln_land_158_lpi_1_dfm_1 | ln_land_159_lpi_1_dfm_1
          | ln_land_163_lpi_1_dfm_1 | ln_land_164_lpi_1_dfm_1 | ln_land_165_lpi_1_dfm_1
          | ln_land_167_lpi_1_dfm_1 | ln_land_168_lpi_1_dfm_1 | ln_land_171_lpi_1_dfm_1
          | ln_land_173_lpi_1_dfm_1 | ln_land_176_lpi_1_dfm_1 | ln_land_178_lpi_1_dfm_1
          | ln_land_179_lpi_1_dfm_1 | ln_land_181_lpi_1_dfm_1 | ln_land_183_lpi_1_dfm_1
          | ln_land_184_lpi_1_dfm_1 | ln_land_187_lpi_1_dfm_1 | ln_land_188_lpi_1_dfm_1
          | ln_land_189_lpi_1_dfm_1 | ln_land_199_lpi_1_dfm_1 | ln_land_200_lpi_1_dfm_1
          | ln_land_203_lpi_1_dfm_1 | ln_land_205_lpi_1_dfm_1 | ln_land_207_lpi_1_dfm_1
          | ln_land_209_lpi_1_dfm_1 | ln_land_210_lpi_1_dfm_1 | ln_land_213_lpi_1_dfm_1
          | ln_land_214_lpi_1_dfm_1 | ln_land_215_lpi_1_dfm_1 | ln_land_216_lpi_1_dfm_1
          | ln_land_217_lpi_1_dfm_1 | ln_land_220_lpi_1_dfm_1 | ln_land_221_lpi_1_dfm_1
          | ln_land_223_lpi_1_dfm_1 | ln_land_224_lpi_1_dfm_1 | ln_land_227_lpi_1_dfm_1
          | ln_land_228_lpi_1_dfm_1 | ln_land_229_lpi_1_dfm_1 | ln_land_232_lpi_1_dfm_1
          | ln_land_234_lpi_1_dfm_1 | ln_land_235_lpi_1_dfm_1 | ln_land_236_lpi_1_dfm_1
          | ln_land_237_lpi_1_dfm_1 | ln_land_238_lpi_1_dfm_1 | ln_land_240_lpi_1_dfm_1)))
          | ln_land_147_lpi_1_dfm_1 | ln_land_148_lpi_1_dfm_1 | ln_land_149_lpi_1_dfm_1
          | ln_land_150_lpi_1_dfm_1 | ln_land_151_lpi_1_dfm_1 | ln_land_152_lpi_1_dfm_1
          | ln_land_153_lpi_1_dfm_1 | ln_land_154_lpi_1_dfm_1 | ln_land_155_lpi_1_dfm_1
          | ln_land_160_lpi_1_dfm_1 | ln_land_161_lpi_1_dfm_1 | ln_land_162_lpi_1_dfm_1
          | ln_land_166_lpi_1_dfm_1 | ln_land_169_lpi_1_dfm_1 | ln_land_170_lpi_1_dfm_1
          | ln_land_172_lpi_1_dfm_1 | ln_land_174_lpi_1_dfm_1 | ln_land_175_lpi_1_dfm_1
          | ln_land_177_lpi_1_dfm_1 | ln_land_180_lpi_1_dfm_1 | ln_land_182_lpi_1_dfm_1
          | ln_land_185_lpi_1_dfm_1 | ln_land_186_lpi_1_dfm_1 | ln_land_190_lpi_1_dfm_1
          | ln_land_191_lpi_1_dfm_1 | ln_land_192_lpi_1_dfm_1 | ln_land_193_lpi_1_dfm_1
          | ln_land_194_lpi_1_dfm_1 | ln_land_195_lpi_1_dfm_1 | ln_land_196_lpi_1_dfm_1
          | ln_land_197_lpi_1_dfm_1 | ln_land_198_lpi_1_dfm_1 | ln_land_201_lpi_1_dfm_1
          | ln_land_202_lpi_1_dfm_1 | ln_land_204_lpi_1_dfm_1 | ln_land_206_lpi_1_dfm_1
          | ln_land_208_lpi_1_dfm_1 | ln_land_211_lpi_1_dfm_1 | ln_land_212_lpi_1_dfm_1
          | ln_land_218_lpi_1_dfm_1 | ln_land_219_lpi_1_dfm_1 | ln_land_222_lpi_1_dfm_1
          | ln_land_225_lpi_1_dfm_1 | ln_land_226_lpi_1_dfm_1 | ln_land_230_lpi_1_dfm_1
          | ln_land_231_lpi_1_dfm_1 | ln_land_233_lpi_1_dfm_1 | ln_land_239_lpi_1_dfm_1
          | ln_land_241_lpi_1_dfm_1 | ln_land_242_lpi_1_dfm_1 | ln_land_243_lpi_1_dfm_1
          | ln_land_244_lpi_1_dfm_1;
      ln_ln_mux1h_118_psp_1_1 <= (((~((~((~((~((((~(((ln_land_4_lpi_1_dfm_1 | ln_and_2_ssc_1
          | ln_land_6_lpi_1_dfm_1) & (~(ln_land_8_lpi_1_dfm_1 | ln_land_9_lpi_1_dfm_1
          | ln_land_10_lpi_1_dfm_1 | ln_land_13_lpi_1_dfm_1 | ln_land_14_lpi_1_dfm_1
          | ln_land_17_lpi_1_dfm_1 | ln_land_19_lpi_1_dfm_1 | ln_land_20_lpi_1_dfm_1
          | ln_land_22_lpi_1_dfm_1 | ln_land_24_lpi_1_dfm_1 | ln_land_26_lpi_1_dfm_1
          | ln_land_29_lpi_1_dfm_1 | ln_land_31_lpi_1_dfm_1 | ln_land_32_lpi_1_dfm_1
          | ln_land_35_lpi_1_dfm_1 | ln_land_36_lpi_1_dfm_1 | ln_land_37_lpi_1_dfm_1
          | ln_land_47_lpi_1_dfm_1 | ln_land_48_lpi_1_dfm_1))) | ln_and_4_ssc_1 |
          ln_land_11_lpi_1_dfm_1 | ln_land_12_lpi_1_dfm_1 | ln_land_15_lpi_1_dfm_1
          | ln_land_16_lpi_1_dfm_1 | ln_land_18_lpi_1_dfm_1 | ln_land_21_lpi_1_dfm_1
          | ln_land_23_lpi_1_dfm_1 | ln_land_25_lpi_1_dfm_1 | ln_land_27_lpi_1_dfm_1
          | ln_land_28_lpi_1_dfm_1 | ln_land_30_lpi_1_dfm_1 | ln_land_33_lpi_1_dfm_1
          | ln_land_34_lpi_1_dfm_1 | ln_land_38_lpi_1_dfm_1 | ln_land_39_lpi_1_dfm_1
          | ln_land_40_lpi_1_dfm_1 | ln_land_41_lpi_1_dfm_1 | ln_land_42_lpi_1_dfm_1
          | ln_land_43_lpi_1_dfm_1 | ln_land_44_lpi_1_dfm_1 | ln_land_45_lpi_1_dfm_1
          | ln_land_46_lpi_1_dfm_1 | ln_land_49_lpi_1_dfm_1 | ln_if_50_ln_if_50_and_seb_1))
          | ln_land_51_lpi_1_dfm_1 | ln_land_52_lpi_1_dfm_1) & (~(ln_and_48_ssc_1
          | ln_land_55_lpi_1_dfm_1 | ln_land_57_lpi_1_dfm_1 | ln_land_59_lpi_1_dfm_1
          | ln_land_62_lpi_1_dfm_1 | ln_land_63_lpi_1_dfm_1 | ln_land_72_lpi_1_dfm_1
          | ln_land_73_lpi_1_dfm_1 | ln_land_75_lpi_1_dfm_1 | ln_land_76_lpi_1_dfm_1
          | ln_land_78_lpi_1_dfm_1 | ln_land_79_lpi_1_dfm_1 | ln_land_81_lpi_1_dfm_1
          | ln_land_82_lpi_1_dfm_1 | ln_land_83_lpi_1_dfm_1 | ln_land_84_lpi_1_dfm_1
          | ln_land_85_lpi_1_dfm_1 | ln_land_86_lpi_1_dfm_1 | ln_land_87_lpi_1_dfm_1
          | ln_land_88_lpi_1_dfm_1 | ln_land_90_lpi_1_dfm_1 | ln_land_92_lpi_1_dfm_1
          | ln_land_94_lpi_1_dfm_1 | ln_land_95_lpi_1_dfm_1 | ln_land_96_lpi_1_dfm_1
          | ln_land_97_lpi_1_dfm_1 | ln_land_98_lpi_1_dfm_1 | ln_land_99_lpi_1_dfm_1
          | ln_land_102_lpi_1_dfm_1 | ln_land_106_lpi_1_dfm_1 | ln_land_109_lpi_1_dfm_1
          | ln_land_111_lpi_1_dfm_1 | ln_land_115_lpi_1_dfm_1 | ln_land_117_lpi_1_dfm_1
          | ln_land_120_lpi_1_dfm_1 | ln_land_121_lpi_1_dfm_1 | ln_land_124_lpi_1_dfm_1
          | ln_land_125_lpi_1_dfm_1 | ln_land_127_lpi_1_dfm_1 | ln_land_130_lpi_1_dfm_1
          | ln_land_132_lpi_1_dfm_1 | ln_land_134_lpi_1_dfm_1 | ln_land_136_lpi_1_dfm_1
          | ln_land_137_lpi_1_dfm_1 | ln_land_139_lpi_1_dfm_1))) | ln_land_54_lpi_1_dfm_1
          | ln_land_56_lpi_1_dfm_1 | ln_land_58_lpi_1_dfm_1 | ln_land_60_lpi_1_dfm_1
          | ln_land_61_lpi_1_dfm_1 | ln_land_64_lpi_1_dfm_1 | ln_land_65_lpi_1_dfm_1
          | ln_land_66_lpi_1_dfm_1 | ln_land_67_lpi_1_dfm_1 | ln_land_68_lpi_1_dfm_1
          | ln_land_69_lpi_1_dfm_1 | ln_land_70_lpi_1_dfm_1 | ln_land_71_lpi_1_dfm_1
          | ln_land_74_lpi_1_dfm_1 | ln_land_77_lpi_1_dfm_1 | ln_land_80_lpi_1_dfm_1
          | ln_land_89_lpi_1_dfm_1 | ln_land_91_lpi_1_dfm_1 | ln_land_93_lpi_1_dfm_1
          | ln_land_100_lpi_1_dfm_1 | ln_land_101_lpi_1_dfm_1 | ln_land_103_lpi_1_dfm_1
          | ln_land_104_lpi_1_dfm_1 | ln_land_105_lpi_1_dfm_1 | ln_land_107_lpi_1_dfm_1
          | ln_land_108_lpi_1_dfm_1 | ln_land_110_lpi_1_dfm_1 | ln_land_112_lpi_1_dfm_1
          | ln_land_113_lpi_1_dfm_1 | ln_land_114_lpi_1_dfm_1 | ln_land_116_lpi_1_dfm_1
          | ln_land_118_lpi_1_dfm_1 | ln_land_119_lpi_1_dfm_1 | ln_land_122_lpi_1_dfm_1
          | ln_land_123_lpi_1_dfm_1 | ln_land_126_lpi_1_dfm_1 | ln_land_128_lpi_1_dfm_1
          | ln_land_129_lpi_1_dfm_1 | ln_land_131_lpi_1_dfm_1 | ln_land_133_lpi_1_dfm_1
          | ln_land_135_lpi_1_dfm_1 | ln_land_138_lpi_1_dfm_1 | ln_land_140_lpi_1_dfm_1))
          | ln_land_142_lpi_1_dfm_1)) | ln_land_141_lpi_1_dfm_1)) | ln_and_138_ssc_1))
          | ln_land_144_lpi_1_dfm_1) & (~(ln_land_147_lpi_1_dfm_1 | ln_land_148_lpi_1_dfm_1
          | ln_land_149_lpi_1_dfm_1 | ln_land_150_lpi_1_dfm_1 | ln_land_151_lpi_1_dfm_1
          | ln_land_152_lpi_1_dfm_1 | ln_land_153_lpi_1_dfm_1 | ln_land_154_lpi_1_dfm_1
          | ln_land_155_lpi_1_dfm_1 | ln_land_159_lpi_1_dfm_1 | ln_land_162_lpi_1_dfm_1
          | ln_land_164_lpi_1_dfm_1 | ln_land_165_lpi_1_dfm_1 | ln_land_168_lpi_1_dfm_1
          | ln_land_170_lpi_1_dfm_1 | ln_land_171_lpi_1_dfm_1 | ln_land_175_lpi_1_dfm_1
          | ln_land_176_lpi_1_dfm_1 | ln_land_177_lpi_1_dfm_1 | ln_land_178_lpi_1_dfm_1
          | ln_land_182_lpi_1_dfm_1 | ln_land_183_lpi_1_dfm_1 | ln_land_185_lpi_1_dfm_1
          | ln_land_187_lpi_1_dfm_1 | ln_land_190_lpi_1_dfm_1 | ln_land_191_lpi_1_dfm_1
          | ln_land_197_lpi_1_dfm_1 | ln_land_198_lpi_1_dfm_1 | ln_land_200_lpi_1_dfm_1
          | ln_land_202_lpi_1_dfm_1 | ln_land_203_lpi_1_dfm_1 | ln_land_209_lpi_1_dfm_1
          | ln_land_211_lpi_1_dfm_1 | ln_land_213_lpi_1_dfm_1 | ln_land_214_lpi_1_dfm_1
          | ln_land_215_lpi_1_dfm_1 | ln_land_216_lpi_1_dfm_1 | ln_land_217_lpi_1_dfm_1
          | ln_land_219_lpi_1_dfm_1 | ln_land_221_lpi_1_dfm_1 | ln_land_222_lpi_1_dfm_1
          | ln_land_223_lpi_1_dfm_1 | ln_land_225_lpi_1_dfm_1 | ln_land_227_lpi_1_dfm_1
          | ln_land_228_lpi_1_dfm_1 | ln_land_229_lpi_1_dfm_1 | ln_land_231_lpi_1_dfm_1
          | ln_land_232_lpi_1_dfm_1 | ln_land_233_lpi_1_dfm_1 | ln_land_234_lpi_1_dfm_1
          | ln_land_238_lpi_1_dfm_1 | ln_land_244_lpi_1_dfm_1))) | ln_and_140_ssc_1
          | ln_land_146_lpi_1_dfm_1 | ln_land_156_lpi_1_dfm_1 | ln_land_157_lpi_1_dfm_1
          | ln_land_158_lpi_1_dfm_1 | ln_land_160_lpi_1_dfm_1 | ln_land_161_lpi_1_dfm_1
          | ln_land_163_lpi_1_dfm_1 | ln_land_166_lpi_1_dfm_1 | ln_land_167_lpi_1_dfm_1
          | ln_land_169_lpi_1_dfm_1 | ln_land_172_lpi_1_dfm_1 | ln_land_173_lpi_1_dfm_1
          | ln_land_174_lpi_1_dfm_1 | ln_land_179_lpi_1_dfm_1 | ln_land_180_lpi_1_dfm_1
          | ln_land_181_lpi_1_dfm_1 | ln_land_184_lpi_1_dfm_1 | ln_land_186_lpi_1_dfm_1
          | ln_land_188_lpi_1_dfm_1 | ln_land_189_lpi_1_dfm_1 | ln_land_192_lpi_1_dfm_1
          | ln_land_193_lpi_1_dfm_1 | ln_land_194_lpi_1_dfm_1 | ln_land_195_lpi_1_dfm_1
          | ln_land_196_lpi_1_dfm_1 | ln_land_199_lpi_1_dfm_1 | ln_land_201_lpi_1_dfm_1
          | ln_land_204_lpi_1_dfm_1 | ln_land_205_lpi_1_dfm_1 | ln_land_206_lpi_1_dfm_1
          | ln_land_207_lpi_1_dfm_1 | ln_land_208_lpi_1_dfm_1 | ln_land_210_lpi_1_dfm_1
          | ln_land_212_lpi_1_dfm_1 | ln_land_218_lpi_1_dfm_1 | ln_land_220_lpi_1_dfm_1
          | ln_land_224_lpi_1_dfm_1 | ln_land_226_lpi_1_dfm_1 | ln_land_230_lpi_1_dfm_1
          | ln_land_235_lpi_1_dfm_1 | ln_land_236_lpi_1_dfm_1 | ln_land_237_lpi_1_dfm_1
          | ln_land_239_lpi_1_dfm_1 | ln_land_240_lpi_1_dfm_1 | ln_land_241_lpi_1_dfm_1
          | ln_land_242_lpi_1_dfm_1 | ln_land_243_lpi_1_dfm_1;
      ln_ln_mux1h_118_psp_1_0 <= (((~((~((~((~((((~((ln_nor_1_cse_1 & (~(ln_land_8_lpi_1_dfm_1
          | ln_land_9_lpi_1_dfm_1 | ln_land_11_lpi_1_dfm_1 | ln_land_13_lpi_1_dfm_1
          | ln_land_15_lpi_1_dfm_1 | ln_land_18_lpi_1_dfm_1 | ln_land_19_lpi_1_dfm_1
          | ln_land_28_lpi_1_dfm_1 | ln_land_29_lpi_1_dfm_1 | ln_land_32_lpi_1_dfm_1
          | ln_land_34_lpi_1_dfm_1 | ln_land_37_lpi_1_dfm_1 | ln_land_41_lpi_1_dfm_1
          | ln_land_42_lpi_1_dfm_1 | ln_land_43_lpi_1_dfm_1 | ln_land_47_lpi_1_dfm_1
          | ln_land_49_lpi_1_dfm_1))) | ln_and_4_ssc_1 | ln_land_10_lpi_1_dfm_1 |
          ln_land_12_lpi_1_dfm_1 | ln_land_14_lpi_1_dfm_1 | ln_land_16_lpi_1_dfm_1
          | ln_land_17_lpi_1_dfm_1 | ln_land_20_lpi_1_dfm_1 | ln_land_21_lpi_1_dfm_1
          | ln_land_22_lpi_1_dfm_1 | ln_land_23_lpi_1_dfm_1 | ln_land_24_lpi_1_dfm_1
          | ln_land_25_lpi_1_dfm_1 | ln_land_26_lpi_1_dfm_1 | ln_land_27_lpi_1_dfm_1
          | ln_land_30_lpi_1_dfm_1 | ln_land_31_lpi_1_dfm_1 | ln_land_33_lpi_1_dfm_1
          | ln_land_35_lpi_1_dfm_1 | ln_land_36_lpi_1_dfm_1 | ln_land_38_lpi_1_dfm_1
          | ln_land_39_lpi_1_dfm_1 | ln_land_40_lpi_1_dfm_1 | ln_land_44_lpi_1_dfm_1
          | ln_land_45_lpi_1_dfm_1 | ln_land_46_lpi_1_dfm_1 | ln_land_48_lpi_1_dfm_1
          | ln_if_50_ln_if_50_and_seb_1 | ln_land_52_lpi_1_dfm_1)) | ln_land_51_lpi_1_dfm_1)
          & (~(ln_and_48_ssc_1 | ln_land_60_lpi_1_dfm_1 | ln_land_62_lpi_1_dfm_1
          | ln_land_64_lpi_1_dfm_1 | ln_land_71_lpi_1_dfm_1 | ln_land_73_lpi_1_dfm_1
          | ln_land_76_lpi_1_dfm_1 | ln_land_77_lpi_1_dfm_1 | ln_land_78_lpi_1_dfm_1
          | ln_land_81_lpi_1_dfm_1 | ln_land_88_lpi_1_dfm_1 | ln_land_94_lpi_1_dfm_1
          | ln_land_99_lpi_1_dfm_1 | ln_land_101_lpi_1_dfm_1 | ln_land_102_lpi_1_dfm_1
          | ln_land_103_lpi_1_dfm_1 | ln_land_106_lpi_1_dfm_1 | ln_land_108_lpi_1_dfm_1
          | ln_land_112_lpi_1_dfm_1 | ln_land_113_lpi_1_dfm_1 | ln_land_114_lpi_1_dfm_1
          | ln_land_118_lpi_1_dfm_1 | ln_land_119_lpi_1_dfm_1 | ln_land_121_lpi_1_dfm_1
          | ln_land_123_lpi_1_dfm_1 | ln_land_125_lpi_1_dfm_1 | ln_land_126_lpi_1_dfm_1
          | ln_land_129_lpi_1_dfm_1 | ln_land_130_lpi_1_dfm_1 | ln_land_131_lpi_1_dfm_1
          | ln_land_132_lpi_1_dfm_1 | ln_land_133_lpi_1_dfm_1 | ln_land_134_lpi_1_dfm_1
          | ln_land_135_lpi_1_dfm_1 | ln_land_136_lpi_1_dfm_1 | ln_land_139_lpi_1_dfm_1
          | ln_land_140_lpi_1_dfm_1))) | ln_land_54_lpi_1_dfm_1 | ln_land_55_lpi_1_dfm_1
          | ln_land_56_lpi_1_dfm_1 | ln_land_57_lpi_1_dfm_1 | ln_land_58_lpi_1_dfm_1
          | ln_land_59_lpi_1_dfm_1 | ln_land_61_lpi_1_dfm_1 | ln_land_63_lpi_1_dfm_1
          | ln_land_65_lpi_1_dfm_1 | ln_land_66_lpi_1_dfm_1 | ln_land_67_lpi_1_dfm_1
          | ln_land_68_lpi_1_dfm_1 | ln_land_69_lpi_1_dfm_1 | ln_land_70_lpi_1_dfm_1
          | ln_land_72_lpi_1_dfm_1 | ln_land_74_lpi_1_dfm_1 | ln_land_75_lpi_1_dfm_1
          | ln_land_79_lpi_1_dfm_1 | ln_land_80_lpi_1_dfm_1 | ln_land_82_lpi_1_dfm_1
          | ln_land_83_lpi_1_dfm_1 | ln_land_84_lpi_1_dfm_1 | ln_land_85_lpi_1_dfm_1
          | ln_land_86_lpi_1_dfm_1 | ln_land_87_lpi_1_dfm_1 | ln_land_89_lpi_1_dfm_1
          | ln_land_90_lpi_1_dfm_1 | ln_land_91_lpi_1_dfm_1 | ln_land_92_lpi_1_dfm_1
          | ln_land_93_lpi_1_dfm_1 | ln_land_95_lpi_1_dfm_1 | ln_land_96_lpi_1_dfm_1
          | ln_land_97_lpi_1_dfm_1 | ln_land_98_lpi_1_dfm_1 | ln_land_100_lpi_1_dfm_1
          | ln_land_104_lpi_1_dfm_1 | ln_land_105_lpi_1_dfm_1 | ln_land_107_lpi_1_dfm_1
          | ln_land_109_lpi_1_dfm_1 | ln_land_110_lpi_1_dfm_1 | ln_land_111_lpi_1_dfm_1
          | ln_land_115_lpi_1_dfm_1 | ln_land_116_lpi_1_dfm_1 | ln_land_117_lpi_1_dfm_1
          | ln_land_120_lpi_1_dfm_1 | ln_land_122_lpi_1_dfm_1 | ln_land_124_lpi_1_dfm_1
          | ln_land_127_lpi_1_dfm_1 | ln_land_128_lpi_1_dfm_1 | ln_land_137_lpi_1_dfm_1
          | ln_land_138_lpi_1_dfm_1)) | ln_land_142_lpi_1_dfm_1)) | ln_land_141_lpi_1_dfm_1))
          | ln_land_144_lpi_1_dfm_1)) | ln_and_138_ssc_1) & (~(ln_land_147_lpi_1_dfm_1
          | ln_land_148_lpi_1_dfm_1 | ln_land_154_lpi_1_dfm_1 | ln_land_155_lpi_1_dfm_1
          | ln_land_157_lpi_1_dfm_1 | ln_land_158_lpi_1_dfm_1 | ln_land_161_lpi_1_dfm_1
          | ln_land_165_lpi_1_dfm_1 | ln_land_166_lpi_1_dfm_1 | ln_land_169_lpi_1_dfm_1
          | ln_land_170_lpi_1_dfm_1 | ln_land_172_lpi_1_dfm_1 | ln_land_175_lpi_1_dfm_1
          | ln_land_176_lpi_1_dfm_1 | ln_land_177_lpi_1_dfm_1 | ln_land_178_lpi_1_dfm_1
          | ln_land_181_lpi_1_dfm_1 | ln_land_183_lpi_1_dfm_1 | ln_land_184_lpi_1_dfm_1
          | ln_land_187_lpi_1_dfm_1 | ln_land_188_lpi_1_dfm_1 | ln_land_192_lpi_1_dfm_1
          | ln_land_193_lpi_1_dfm_1 | ln_land_194_lpi_1_dfm_1 | ln_land_195_lpi_1_dfm_1
          | ln_land_196_lpi_1_dfm_1 | ln_land_198_lpi_1_dfm_1 | ln_land_199_lpi_1_dfm_1
          | ln_land_200_lpi_1_dfm_1 | ln_land_201_lpi_1_dfm_1 | ln_land_202_lpi_1_dfm_1
          | ln_land_204_lpi_1_dfm_1 | ln_land_207_lpi_1_dfm_1 | ln_land_208_lpi_1_dfm_1
          | ln_land_213_lpi_1_dfm_1 | ln_land_217_lpi_1_dfm_1 | ln_land_221_lpi_1_dfm_1
          | ln_land_222_lpi_1_dfm_1 | ln_land_223_lpi_1_dfm_1 | ln_land_227_lpi_1_dfm_1
          | ln_land_228_lpi_1_dfm_1 | ln_land_229_lpi_1_dfm_1 | ln_land_230_lpi_1_dfm_1
          | ln_land_231_lpi_1_dfm_1 | ln_land_234_lpi_1_dfm_1 | ln_land_235_lpi_1_dfm_1
          | ln_land_241_lpi_1_dfm_1))) | ln_and_140_ssc_1 | ln_land_146_lpi_1_dfm_1
          | ln_land_149_lpi_1_dfm_1 | ln_land_150_lpi_1_dfm_1 | ln_land_151_lpi_1_dfm_1
          | ln_land_152_lpi_1_dfm_1 | ln_land_153_lpi_1_dfm_1 | ln_land_156_lpi_1_dfm_1
          | ln_land_159_lpi_1_dfm_1 | ln_land_160_lpi_1_dfm_1 | ln_land_162_lpi_1_dfm_1
          | ln_land_163_lpi_1_dfm_1 | ln_land_164_lpi_1_dfm_1 | ln_land_167_lpi_1_dfm_1
          | ln_land_168_lpi_1_dfm_1 | ln_land_171_lpi_1_dfm_1 | ln_land_173_lpi_1_dfm_1
          | ln_land_174_lpi_1_dfm_1 | ln_land_179_lpi_1_dfm_1 | ln_land_180_lpi_1_dfm_1
          | ln_land_182_lpi_1_dfm_1 | ln_land_185_lpi_1_dfm_1 | ln_land_186_lpi_1_dfm_1
          | ln_land_189_lpi_1_dfm_1 | ln_land_190_lpi_1_dfm_1 | ln_land_191_lpi_1_dfm_1
          | ln_land_197_lpi_1_dfm_1 | ln_land_203_lpi_1_dfm_1 | ln_land_205_lpi_1_dfm_1
          | ln_land_206_lpi_1_dfm_1 | ln_land_209_lpi_1_dfm_1 | ln_land_210_lpi_1_dfm_1
          | ln_land_211_lpi_1_dfm_1 | ln_land_212_lpi_1_dfm_1 | ln_land_214_lpi_1_dfm_1
          | ln_land_215_lpi_1_dfm_1 | ln_land_216_lpi_1_dfm_1 | ln_land_218_lpi_1_dfm_1
          | ln_land_219_lpi_1_dfm_1 | ln_land_220_lpi_1_dfm_1 | ln_land_224_lpi_1_dfm_1
          | ln_land_225_lpi_1_dfm_1 | ln_land_226_lpi_1_dfm_1 | ln_land_232_lpi_1_dfm_1
          | ln_land_233_lpi_1_dfm_1 | ln_land_236_lpi_1_dfm_1 | ln_land_237_lpi_1_dfm_1
          | ln_land_238_lpi_1_dfm_1 | ln_land_239_lpi_1_dfm_1 | ln_land_240_lpi_1_dfm_1
          | ln_land_242_lpi_1_dfm_1 | ln_land_243_lpi_1_dfm_1 | ln_land_244_lpi_1_dfm_1;
      operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1 <= operator_24_14_false_AC_TRN_AC_WRAP_slc_P1_24_23_0_cse_23_10_sva_1_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      sum2_1_lpi_1_dfm_1 <= 24'b000000000000000000000000;
    end
    else if ( MUX_s_1_2_2(and_277_nl, and_276_cse, or_2_tmp) ) begin
      sum2_1_lpi_1_dfm_1 <= MUX_v_24_2_2(24'b000000000000000000000000, sum2_1_lpi_1_dfm_1_mx0,
          if_4_for_if_4_for_if_4_for_not_2_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      ln_1_land_251_lpi_1_dfm_1 <= 1'b0;
      ln_1_land_252_lpi_1_dfm_1 <= 1'b0;
      ln_1_ln_1_mux1h_118_psp_1_12 <= 1'b0;
      ln_1_and_248_ssc_1 <= 1'b0;
      ln_1_if_253_acc_cse_11_sva_1 <= 1'b0;
      ln_1_ln_1_mux1h_118_psp_1_11 <= 1'b0;
      ln_1_ln_1_mux1h_118_psp_1_10 <= 1'b0;
      ln_1_and_407_ssc_1 <= 1'b0;
      ln_1_and_244_ssc_1 <= 1'b0;
      ln_1_and_379_ssc_1 <= 1'b0;
      ln_1_and_240_ssc_1 <= 1'b0;
      ln_1_and_377_ssc_1 <= 1'b0;
      ln_1_and_242_ssc_1 <= 1'b0;
      ln_1_and_427_itm_1 <= 1'b0;
      ln_1_ln_1_mux1h_118_psp_1_8 <= 1'b0;
      ln_1_ln_1_mux1h_118_psp_1_7 <= 1'b0;
      ln_1_ln_1_mux1h_118_psp_1_6 <= 1'b0;
      ln_1_ln_1_mux1h_118_psp_1_5 <= 1'b0;
      ln_1_ln_1_mux1h_118_psp_1_4 <= 1'b0;
      ln_1_ln_1_mux1h_118_psp_1_3 <= 1'b0;
      ln_1_ln_1_mux1h_118_psp_1_2 <= 1'b0;
      ln_1_ln_1_mux1h_118_psp_1_1 <= 1'b0;
      ln_1_ln_1_mux1h_118_psp_1_0 <= 1'b0;
      operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1
          <= 14'b00000000000000;
    end
    else if ( and_dcpl_61 ) begin
      ln_1_land_251_lpi_1_dfm_1 <= ln_1_land_251_lpi_1_dfm_1_1;
      ln_1_land_252_lpi_1_dfm_1 <= ln_1_land_252_lpi_1_dfm_1_1;
      ln_1_ln_1_mux1h_118_psp_1_12 <= (~(ln_1_land_141_lpi_1_dfm_1 | ln_1_land_142_lpi_1_dfm_1))
          & ln_1_nor_3_cse_1 & (~(ln_1_and_140_ssc_1 | ln_1_land_146_lpi_1_dfm_1
          | ln_1_land_147_lpi_1_dfm_1 | ln_1_land_148_lpi_1_dfm_1 | ln_1_land_149_lpi_1_dfm_1
          | ln_1_land_150_lpi_1_dfm_1 | ln_1_land_151_lpi_1_dfm_1 | ln_1_land_152_lpi_1_dfm_1
          | ln_1_land_153_lpi_1_dfm_1 | ln_1_land_154_lpi_1_dfm_1 | ln_1_land_155_lpi_1_dfm_1
          | ln_1_land_156_lpi_1_dfm_1 | ln_1_land_157_lpi_1_dfm_1 | ln_1_land_158_lpi_1_dfm_1
          | ln_1_land_159_lpi_1_dfm_1 | ln_1_land_160_lpi_1_dfm_1 | ln_1_land_161_lpi_1_dfm_1
          | ln_1_land_162_lpi_1_dfm_1 | ln_1_land_163_lpi_1_dfm_1 | ln_1_land_164_lpi_1_dfm_1
          | ln_1_land_165_lpi_1_dfm_1 | ln_1_land_166_lpi_1_dfm_1 | ln_1_land_167_lpi_1_dfm_1
          | ln_1_land_168_lpi_1_dfm_1 | ln_1_land_169_lpi_1_dfm_1 | ln_1_land_170_lpi_1_dfm_1
          | ln_1_land_171_lpi_1_dfm_1 | ln_1_land_172_lpi_1_dfm_1 | ln_1_land_173_lpi_1_dfm_1
          | ln_1_land_174_lpi_1_dfm_1 | ln_1_land_175_lpi_1_dfm_1 | ln_1_land_176_lpi_1_dfm_1
          | ln_1_land_177_lpi_1_dfm_1 | ln_1_land_178_lpi_1_dfm_1 | ln_1_land_179_lpi_1_dfm_1
          | ln_1_land_180_lpi_1_dfm_1 | ln_1_land_181_lpi_1_dfm_1 | ln_1_land_182_lpi_1_dfm_1
          | ln_1_land_183_lpi_1_dfm_1 | ln_1_land_184_lpi_1_dfm_1 | ln_1_land_185_lpi_1_dfm_1
          | ln_1_land_186_lpi_1_dfm_1 | ln_1_land_187_lpi_1_dfm_1 | ln_1_land_188_lpi_1_dfm_1
          | ln_1_land_189_lpi_1_dfm_1 | ln_1_land_190_lpi_1_dfm_1 | ln_1_land_191_lpi_1_dfm_1
          | ln_1_land_192_lpi_1_dfm_1 | ln_1_land_193_lpi_1_dfm_1 | ln_1_land_194_lpi_1_dfm_1
          | ln_1_land_195_lpi_1_dfm_1 | ln_1_land_196_lpi_1_dfm_1 | ln_1_land_197_lpi_1_dfm_1
          | ln_1_land_198_lpi_1_dfm_1 | ln_1_land_199_lpi_1_dfm_1 | ln_1_land_200_lpi_1_dfm_1
          | ln_1_land_201_lpi_1_dfm_1 | ln_1_land_202_lpi_1_dfm_1 | ln_1_land_203_lpi_1_dfm_1
          | ln_1_land_204_lpi_1_dfm_1 | ln_1_land_205_lpi_1_dfm_1 | ln_1_land_206_lpi_1_dfm_1
          | ln_1_land_207_lpi_1_dfm_1 | ln_1_land_208_lpi_1_dfm_1 | ln_1_land_209_lpi_1_dfm_1
          | ln_1_land_210_lpi_1_dfm_1 | ln_1_land_211_lpi_1_dfm_1 | ln_1_land_212_lpi_1_dfm_1
          | ln_1_land_213_lpi_1_dfm_1 | ln_1_land_214_lpi_1_dfm_1 | ln_1_land_215_lpi_1_dfm_1
          | ln_1_land_216_lpi_1_dfm_1 | ln_1_land_217_lpi_1_dfm_1 | ln_1_land_218_lpi_1_dfm_1
          | ln_1_land_219_lpi_1_dfm_1 | ln_1_land_220_lpi_1_dfm_1 | ln_1_land_221_lpi_1_dfm_1
          | ln_1_land_222_lpi_1_dfm_1 | ln_1_land_223_lpi_1_dfm_1 | ln_1_land_224_lpi_1_dfm_1
          | ln_1_land_225_lpi_1_dfm_1 | ln_1_land_226_lpi_1_dfm_1 | ln_1_land_227_lpi_1_dfm_1
          | ln_1_land_228_lpi_1_dfm_1 | ln_1_land_229_lpi_1_dfm_1 | ln_1_land_230_lpi_1_dfm_1
          | ln_1_land_231_lpi_1_dfm_1 | ln_1_land_232_lpi_1_dfm_1 | ln_1_land_233_lpi_1_dfm_1
          | ln_1_land_234_lpi_1_dfm_1 | ln_1_land_235_lpi_1_dfm_1 | ln_1_land_236_lpi_1_dfm_1
          | ln_1_land_237_lpi_1_dfm_1 | ln_1_land_238_lpi_1_dfm_1 | ln_1_land_239_lpi_1_dfm_1
          | ln_1_land_240_lpi_1_dfm_1 | ln_1_land_241_lpi_1_dfm_1 | ln_1_land_242_lpi_1_dfm_1
          | ln_1_land_243_lpi_1_dfm_1 | ln_1_land_244_lpi_1_dfm_1));
      ln_1_and_248_ssc_1 <= ln_1_if_252_acc_itm_12_1 & (~ ln_1_if_253_acc_itm_11_1);
      ln_1_if_253_acc_cse_11_sva_1 <= ln_1_if_253_acc_itm_11_1;
      ln_1_ln_1_mux1h_118_psp_1_11 <= ((((~(ln_1_land_51_lpi_1_dfm_1 | ln_1_land_52_lpi_1_dfm_1))
          & (~(ln_1_and_48_ssc_1 | ln_1_land_54_lpi_1_dfm_1 | ln_1_land_55_lpi_1_dfm_1
          | ln_1_land_56_lpi_1_dfm_1 | ln_1_land_57_lpi_1_dfm_1 | ln_1_land_58_lpi_1_dfm_1
          | ln_1_land_59_lpi_1_dfm_1 | ln_1_land_60_lpi_1_dfm_1 | ln_1_land_61_lpi_1_dfm_1
          | ln_1_land_62_lpi_1_dfm_1 | ln_1_land_63_lpi_1_dfm_1 | ln_1_land_64_lpi_1_dfm_1
          | ln_1_land_65_lpi_1_dfm_1 | ln_1_land_66_lpi_1_dfm_1 | ln_1_land_67_lpi_1_dfm_1
          | ln_1_land_68_lpi_1_dfm_1 | ln_1_land_69_lpi_1_dfm_1 | ln_1_land_70_lpi_1_dfm_1
          | ln_1_land_71_lpi_1_dfm_1 | ln_1_land_72_lpi_1_dfm_1 | ln_1_land_73_lpi_1_dfm_1
          | ln_1_land_74_lpi_1_dfm_1 | ln_1_land_75_lpi_1_dfm_1 | ln_1_land_76_lpi_1_dfm_1
          | ln_1_land_77_lpi_1_dfm_1 | ln_1_land_78_lpi_1_dfm_1 | ln_1_land_79_lpi_1_dfm_1
          | ln_1_land_80_lpi_1_dfm_1 | ln_1_land_81_lpi_1_dfm_1 | ln_1_land_82_lpi_1_dfm_1
          | ln_1_land_83_lpi_1_dfm_1 | ln_1_land_84_lpi_1_dfm_1 | ln_1_land_85_lpi_1_dfm_1
          | ln_1_land_86_lpi_1_dfm_1 | ln_1_land_87_lpi_1_dfm_1 | ln_1_land_88_lpi_1_dfm_1
          | ln_1_land_89_lpi_1_dfm_1 | ln_1_land_90_lpi_1_dfm_1 | ln_1_land_91_lpi_1_dfm_1
          | ln_1_land_92_lpi_1_dfm_1 | ln_1_land_93_lpi_1_dfm_1 | ln_1_land_94_lpi_1_dfm_1
          | ln_1_land_95_lpi_1_dfm_1 | ln_1_land_96_lpi_1_dfm_1 | ln_1_land_97_lpi_1_dfm_1
          | ln_1_land_98_lpi_1_dfm_1 | ln_1_land_99_lpi_1_dfm_1 | ln_1_land_100_lpi_1_dfm_1
          | ln_1_land_101_lpi_1_dfm_1 | ln_1_land_102_lpi_1_dfm_1 | ln_1_land_103_lpi_1_dfm_1
          | ln_1_land_104_lpi_1_dfm_1 | ln_1_land_105_lpi_1_dfm_1 | ln_1_land_106_lpi_1_dfm_1
          | ln_1_land_107_lpi_1_dfm_1 | ln_1_land_108_lpi_1_dfm_1 | ln_1_land_109_lpi_1_dfm_1
          | ln_1_land_110_lpi_1_dfm_1 | ln_1_land_111_lpi_1_dfm_1 | ln_1_land_112_lpi_1_dfm_1
          | ln_1_land_113_lpi_1_dfm_1 | ln_1_land_114_lpi_1_dfm_1 | ln_1_land_115_lpi_1_dfm_1
          | ln_1_land_116_lpi_1_dfm_1 | ln_1_land_117_lpi_1_dfm_1 | ln_1_land_118_lpi_1_dfm_1
          | ln_1_land_119_lpi_1_dfm_1 | ln_1_land_120_lpi_1_dfm_1 | ln_1_land_121_lpi_1_dfm_1
          | ln_1_land_122_lpi_1_dfm_1 | ln_1_land_123_lpi_1_dfm_1 | ln_1_land_124_lpi_1_dfm_1
          | ln_1_land_125_lpi_1_dfm_1 | ln_1_land_126_lpi_1_dfm_1 | ln_1_land_127_lpi_1_dfm_1
          | ln_1_land_128_lpi_1_dfm_1 | ln_1_land_129_lpi_1_dfm_1 | ln_1_land_130_lpi_1_dfm_1
          | ln_1_land_131_lpi_1_dfm_1 | ln_1_land_132_lpi_1_dfm_1 | ln_1_land_133_lpi_1_dfm_1
          | ln_1_land_134_lpi_1_dfm_1 | ln_1_land_135_lpi_1_dfm_1 | ln_1_land_136_lpi_1_dfm_1
          | ln_1_land_137_lpi_1_dfm_1 | ln_1_land_138_lpi_1_dfm_1 | ln_1_land_139_lpi_1_dfm_1
          | ln_1_land_140_lpi_1_dfm_1))) | ln_1_land_141_lpi_1_dfm_1 | ln_1_land_142_lpi_1_dfm_1
          | ln_1_and_138_ssc_1 | ln_1_land_144_lpi_1_dfm_1) & ln_1_and_368_m1c_1)
          | ln_1_and_140_ssc_1 | ln_1_land_146_lpi_1_dfm_1 | ln_1_land_147_lpi_1_dfm_1
          | ln_1_land_148_lpi_1_dfm_1 | ln_1_land_149_lpi_1_dfm_1 | ln_1_land_150_lpi_1_dfm_1
          | ln_1_land_151_lpi_1_dfm_1 | ln_1_land_152_lpi_1_dfm_1 | ln_1_land_153_lpi_1_dfm_1
          | ln_1_land_154_lpi_1_dfm_1 | ln_1_land_155_lpi_1_dfm_1 | ln_1_land_156_lpi_1_dfm_1
          | ln_1_land_157_lpi_1_dfm_1 | ln_1_land_158_lpi_1_dfm_1 | ln_1_land_159_lpi_1_dfm_1
          | ln_1_land_160_lpi_1_dfm_1 | ln_1_land_161_lpi_1_dfm_1 | ln_1_land_162_lpi_1_dfm_1
          | ln_1_land_163_lpi_1_dfm_1 | ln_1_land_164_lpi_1_dfm_1 | ln_1_land_165_lpi_1_dfm_1
          | ln_1_land_166_lpi_1_dfm_1 | ln_1_land_167_lpi_1_dfm_1 | ln_1_land_168_lpi_1_dfm_1
          | ln_1_land_169_lpi_1_dfm_1 | ln_1_land_170_lpi_1_dfm_1 | ln_1_land_171_lpi_1_dfm_1
          | ln_1_land_172_lpi_1_dfm_1 | ln_1_land_173_lpi_1_dfm_1 | ln_1_land_174_lpi_1_dfm_1
          | ln_1_land_175_lpi_1_dfm_1 | ln_1_land_176_lpi_1_dfm_1 | ln_1_land_177_lpi_1_dfm_1
          | ln_1_land_178_lpi_1_dfm_1 | ln_1_land_179_lpi_1_dfm_1 | ln_1_land_180_lpi_1_dfm_1
          | ln_1_land_181_lpi_1_dfm_1 | ln_1_land_182_lpi_1_dfm_1 | ln_1_land_183_lpi_1_dfm_1
          | ln_1_land_184_lpi_1_dfm_1 | ln_1_land_185_lpi_1_dfm_1 | ln_1_land_186_lpi_1_dfm_1
          | ln_1_land_187_lpi_1_dfm_1 | ln_1_land_188_lpi_1_dfm_1 | ln_1_land_189_lpi_1_dfm_1
          | ln_1_land_190_lpi_1_dfm_1 | ln_1_land_191_lpi_1_dfm_1 | ln_1_land_192_lpi_1_dfm_1
          | ln_1_land_193_lpi_1_dfm_1 | ln_1_land_194_lpi_1_dfm_1 | ln_1_land_195_lpi_1_dfm_1
          | ln_1_land_196_lpi_1_dfm_1 | ln_1_land_197_lpi_1_dfm_1 | ln_1_land_198_lpi_1_dfm_1
          | ln_1_land_199_lpi_1_dfm_1 | ln_1_land_200_lpi_1_dfm_1 | ln_1_land_201_lpi_1_dfm_1
          | ln_1_land_202_lpi_1_dfm_1 | ln_1_land_203_lpi_1_dfm_1 | ln_1_land_204_lpi_1_dfm_1
          | ln_1_land_205_lpi_1_dfm_1 | ln_1_land_206_lpi_1_dfm_1 | ln_1_land_207_lpi_1_dfm_1
          | ln_1_land_208_lpi_1_dfm_1 | ln_1_land_209_lpi_1_dfm_1 | ln_1_land_210_lpi_1_dfm_1
          | ln_1_land_211_lpi_1_dfm_1 | ln_1_land_212_lpi_1_dfm_1 | ln_1_land_213_lpi_1_dfm_1
          | ln_1_land_214_lpi_1_dfm_1 | ln_1_land_215_lpi_1_dfm_1 | ln_1_land_216_lpi_1_dfm_1
          | ln_1_land_217_lpi_1_dfm_1 | ln_1_land_218_lpi_1_dfm_1 | ln_1_land_219_lpi_1_dfm_1
          | ln_1_land_220_lpi_1_dfm_1 | ln_1_land_221_lpi_1_dfm_1 | ln_1_land_222_lpi_1_dfm_1
          | ln_1_land_223_lpi_1_dfm_1 | ln_1_land_224_lpi_1_dfm_1 | ln_1_land_225_lpi_1_dfm_1
          | ln_1_land_226_lpi_1_dfm_1 | ln_1_land_227_lpi_1_dfm_1 | ln_1_land_228_lpi_1_dfm_1;
      ln_1_ln_1_mux1h_118_psp_1_10 <= (((((~(ln_1_land_6_lpi_1_dfm_1 | ln_1_and_4_ssc_1
          | ln_1_land_8_lpi_1_dfm_1 | ln_1_land_9_lpi_1_dfm_1 | ln_1_land_10_lpi_1_dfm_1
          | ln_1_land_11_lpi_1_dfm_1 | ln_1_land_12_lpi_1_dfm_1 | ln_1_land_13_lpi_1_dfm_1
          | ln_1_land_14_lpi_1_dfm_1 | ln_1_land_15_lpi_1_dfm_1 | ln_1_land_16_lpi_1_dfm_1
          | ln_1_land_17_lpi_1_dfm_1 | ln_1_land_18_lpi_1_dfm_1 | ln_1_land_19_lpi_1_dfm_1
          | ln_1_land_20_lpi_1_dfm_1 | ln_1_land_21_lpi_1_dfm_1 | ln_1_land_22_lpi_1_dfm_1
          | ln_1_land_23_lpi_1_dfm_1 | ln_1_land_24_lpi_1_dfm_1 | ln_1_land_25_lpi_1_dfm_1
          | ln_1_land_26_lpi_1_dfm_1 | ln_1_land_27_lpi_1_dfm_1 | ln_1_land_28_lpi_1_dfm_1
          | ln_1_land_29_lpi_1_dfm_1 | ln_1_land_30_lpi_1_dfm_1 | ln_1_land_31_lpi_1_dfm_1
          | ln_1_land_32_lpi_1_dfm_1 | ln_1_land_33_lpi_1_dfm_1 | ln_1_land_34_lpi_1_dfm_1
          | ln_1_land_35_lpi_1_dfm_1 | ln_1_land_36_lpi_1_dfm_1 | ln_1_land_37_lpi_1_dfm_1
          | ln_1_land_38_lpi_1_dfm_1 | ln_1_land_39_lpi_1_dfm_1 | ln_1_land_40_lpi_1_dfm_1
          | ln_1_land_41_lpi_1_dfm_1 | ln_1_land_42_lpi_1_dfm_1 | ln_1_land_43_lpi_1_dfm_1
          | ln_1_land_44_lpi_1_dfm_1 | ln_1_land_45_lpi_1_dfm_1 | ln_1_land_46_lpi_1_dfm_1
          | ln_1_land_47_lpi_1_dfm_1 | ln_1_land_48_lpi_1_dfm_1 | ln_1_land_49_lpi_1_dfm_1
          | ln_1_if_50_ln_1_if_50_and_seb_1)) | ln_1_land_51_lpi_1_dfm_1 | ln_1_land_52_lpi_1_dfm_1)
          & (~(ln_1_land_98_lpi_1_dfm_1 | ln_1_land_99_lpi_1_dfm_1 | ln_1_land_100_lpi_1_dfm_1
          | ln_1_land_101_lpi_1_dfm_1 | ln_1_land_102_lpi_1_dfm_1 | ln_1_land_103_lpi_1_dfm_1
          | ln_1_land_104_lpi_1_dfm_1 | ln_1_land_105_lpi_1_dfm_1 | ln_1_land_106_lpi_1_dfm_1
          | ln_1_land_107_lpi_1_dfm_1 | ln_1_land_108_lpi_1_dfm_1 | ln_1_land_109_lpi_1_dfm_1
          | ln_1_land_110_lpi_1_dfm_1 | ln_1_land_111_lpi_1_dfm_1 | ln_1_land_112_lpi_1_dfm_1
          | ln_1_land_113_lpi_1_dfm_1 | ln_1_land_114_lpi_1_dfm_1 | ln_1_land_115_lpi_1_dfm_1
          | ln_1_land_116_lpi_1_dfm_1 | ln_1_land_117_lpi_1_dfm_1 | ln_1_land_118_lpi_1_dfm_1
          | ln_1_land_119_lpi_1_dfm_1 | ln_1_land_120_lpi_1_dfm_1 | ln_1_land_121_lpi_1_dfm_1
          | ln_1_land_122_lpi_1_dfm_1 | ln_1_land_123_lpi_1_dfm_1 | ln_1_land_124_lpi_1_dfm_1
          | ln_1_land_125_lpi_1_dfm_1 | ln_1_land_126_lpi_1_dfm_1 | ln_1_land_127_lpi_1_dfm_1
          | ln_1_land_128_lpi_1_dfm_1 | ln_1_land_129_lpi_1_dfm_1 | ln_1_land_130_lpi_1_dfm_1
          | ln_1_land_131_lpi_1_dfm_1 | ln_1_land_132_lpi_1_dfm_1 | ln_1_land_133_lpi_1_dfm_1
          | ln_1_land_134_lpi_1_dfm_1 | ln_1_land_135_lpi_1_dfm_1 | ln_1_land_136_lpi_1_dfm_1
          | ln_1_land_137_lpi_1_dfm_1 | ln_1_land_138_lpi_1_dfm_1 | ln_1_land_139_lpi_1_dfm_1
          | ln_1_land_140_lpi_1_dfm_1))) | ln_1_and_48_ssc_1 | ln_1_land_54_lpi_1_dfm_1
          | ln_1_land_55_lpi_1_dfm_1 | ln_1_land_56_lpi_1_dfm_1 | ln_1_land_57_lpi_1_dfm_1
          | ln_1_land_58_lpi_1_dfm_1 | ln_1_land_59_lpi_1_dfm_1 | ln_1_land_60_lpi_1_dfm_1
          | ln_1_land_61_lpi_1_dfm_1 | ln_1_land_62_lpi_1_dfm_1 | ln_1_land_63_lpi_1_dfm_1
          | ln_1_land_64_lpi_1_dfm_1 | ln_1_land_65_lpi_1_dfm_1 | ln_1_land_66_lpi_1_dfm_1
          | ln_1_land_67_lpi_1_dfm_1 | ln_1_land_68_lpi_1_dfm_1 | ln_1_land_69_lpi_1_dfm_1
          | ln_1_land_70_lpi_1_dfm_1 | ln_1_land_71_lpi_1_dfm_1 | ln_1_land_72_lpi_1_dfm_1
          | ln_1_land_73_lpi_1_dfm_1 | ln_1_land_74_lpi_1_dfm_1 | ln_1_land_75_lpi_1_dfm_1
          | ln_1_land_76_lpi_1_dfm_1 | ln_1_land_77_lpi_1_dfm_1 | ln_1_land_78_lpi_1_dfm_1
          | ln_1_land_79_lpi_1_dfm_1 | ln_1_land_80_lpi_1_dfm_1 | ln_1_land_81_lpi_1_dfm_1
          | ln_1_land_82_lpi_1_dfm_1 | ln_1_land_83_lpi_1_dfm_1 | ln_1_land_84_lpi_1_dfm_1
          | ln_1_land_85_lpi_1_dfm_1 | ln_1_land_86_lpi_1_dfm_1 | ln_1_land_87_lpi_1_dfm_1
          | ln_1_land_88_lpi_1_dfm_1 | ln_1_land_89_lpi_1_dfm_1 | ln_1_land_90_lpi_1_dfm_1
          | ln_1_land_91_lpi_1_dfm_1 | ln_1_land_92_lpi_1_dfm_1 | ln_1_land_93_lpi_1_dfm_1
          | ln_1_land_94_lpi_1_dfm_1 | ln_1_land_95_lpi_1_dfm_1 | ln_1_land_96_lpi_1_dfm_1
          | ln_1_land_97_lpi_1_dfm_1 | ln_1_land_141_lpi_1_dfm_1 | ln_1_land_142_lpi_1_dfm_1
          | ln_1_and_138_ssc_1 | ln_1_land_144_lpi_1_dfm_1) & (~(ln_1_land_195_lpi_1_dfm_1
          | ln_1_land_196_lpi_1_dfm_1 | ln_1_land_197_lpi_1_dfm_1 | ln_1_land_198_lpi_1_dfm_1
          | ln_1_land_199_lpi_1_dfm_1 | ln_1_land_200_lpi_1_dfm_1 | ln_1_land_201_lpi_1_dfm_1
          | ln_1_land_202_lpi_1_dfm_1 | ln_1_land_203_lpi_1_dfm_1 | ln_1_land_204_lpi_1_dfm_1
          | ln_1_land_205_lpi_1_dfm_1 | ln_1_land_206_lpi_1_dfm_1 | ln_1_land_207_lpi_1_dfm_1
          | ln_1_land_208_lpi_1_dfm_1 | ln_1_land_209_lpi_1_dfm_1 | ln_1_land_210_lpi_1_dfm_1
          | ln_1_land_211_lpi_1_dfm_1 | ln_1_land_212_lpi_1_dfm_1 | ln_1_land_213_lpi_1_dfm_1
          | ln_1_land_214_lpi_1_dfm_1 | ln_1_land_215_lpi_1_dfm_1 | ln_1_land_216_lpi_1_dfm_1
          | ln_1_land_217_lpi_1_dfm_1 | ln_1_land_218_lpi_1_dfm_1 | ln_1_land_219_lpi_1_dfm_1
          | ln_1_land_220_lpi_1_dfm_1 | ln_1_land_221_lpi_1_dfm_1 | ln_1_land_222_lpi_1_dfm_1
          | ln_1_land_223_lpi_1_dfm_1 | ln_1_land_224_lpi_1_dfm_1 | ln_1_land_225_lpi_1_dfm_1
          | ln_1_land_226_lpi_1_dfm_1 | ln_1_land_227_lpi_1_dfm_1 | ln_1_land_228_lpi_1_dfm_1)))
          | ln_1_and_140_ssc_1 | ln_1_land_146_lpi_1_dfm_1 | ln_1_land_147_lpi_1_dfm_1
          | ln_1_land_148_lpi_1_dfm_1 | ln_1_land_149_lpi_1_dfm_1 | ln_1_land_150_lpi_1_dfm_1
          | ln_1_land_151_lpi_1_dfm_1 | ln_1_land_152_lpi_1_dfm_1 | ln_1_land_153_lpi_1_dfm_1
          | ln_1_land_154_lpi_1_dfm_1 | ln_1_land_155_lpi_1_dfm_1 | ln_1_land_156_lpi_1_dfm_1
          | ln_1_land_157_lpi_1_dfm_1 | ln_1_land_158_lpi_1_dfm_1 | ln_1_land_159_lpi_1_dfm_1
          | ln_1_land_160_lpi_1_dfm_1 | ln_1_land_161_lpi_1_dfm_1 | ln_1_land_162_lpi_1_dfm_1
          | ln_1_land_163_lpi_1_dfm_1 | ln_1_land_164_lpi_1_dfm_1 | ln_1_land_165_lpi_1_dfm_1
          | ln_1_land_166_lpi_1_dfm_1 | ln_1_land_167_lpi_1_dfm_1 | ln_1_land_168_lpi_1_dfm_1
          | ln_1_land_169_lpi_1_dfm_1 | ln_1_land_170_lpi_1_dfm_1 | ln_1_land_171_lpi_1_dfm_1
          | ln_1_land_172_lpi_1_dfm_1 | ln_1_land_173_lpi_1_dfm_1 | ln_1_land_174_lpi_1_dfm_1
          | ln_1_land_175_lpi_1_dfm_1 | ln_1_land_176_lpi_1_dfm_1 | ln_1_land_177_lpi_1_dfm_1
          | ln_1_land_178_lpi_1_dfm_1 | ln_1_land_179_lpi_1_dfm_1 | ln_1_land_180_lpi_1_dfm_1
          | ln_1_land_181_lpi_1_dfm_1 | ln_1_land_182_lpi_1_dfm_1 | ln_1_land_183_lpi_1_dfm_1
          | ln_1_land_184_lpi_1_dfm_1 | ln_1_land_185_lpi_1_dfm_1 | ln_1_land_186_lpi_1_dfm_1
          | ln_1_land_187_lpi_1_dfm_1 | ln_1_land_188_lpi_1_dfm_1 | ln_1_land_189_lpi_1_dfm_1
          | ln_1_land_190_lpi_1_dfm_1 | ln_1_land_191_lpi_1_dfm_1 | ln_1_land_192_lpi_1_dfm_1
          | ln_1_land_193_lpi_1_dfm_1 | ln_1_land_194_lpi_1_dfm_1 | ln_1_land_229_lpi_1_dfm_1
          | ln_1_land_230_lpi_1_dfm_1 | ln_1_land_231_lpi_1_dfm_1 | ln_1_land_232_lpi_1_dfm_1
          | ln_1_land_233_lpi_1_dfm_1 | ln_1_land_234_lpi_1_dfm_1 | ln_1_land_235_lpi_1_dfm_1
          | ln_1_land_236_lpi_1_dfm_1 | ln_1_land_237_lpi_1_dfm_1 | ln_1_land_238_lpi_1_dfm_1
          | ln_1_land_239_lpi_1_dfm_1 | ln_1_land_240_lpi_1_dfm_1 | ln_1_land_241_lpi_1_dfm_1
          | ln_1_land_242_lpi_1_dfm_1 | ln_1_land_243_lpi_1_dfm_1 | ln_1_land_244_lpi_1_dfm_1;
      ln_1_and_407_ssc_1 <= ln_1_land_248_lpi_1_dfm_1;
      ln_1_and_244_ssc_1 <= ln_1_land_249_lpi_1_dfm_1;
      ln_1_and_379_ssc_1 <= ln_1_land_250_lpi_1_dfm_1;
      ln_1_and_240_ssc_1 <= ln_1_and_240_ssc_1_1;
      ln_1_and_377_ssc_1 <= ln_1_land_246_lpi_1_dfm_1;
      ln_1_and_242_ssc_1 <= ln_1_land_247_lpi_1_dfm_1;
      ln_1_and_427_itm_1 <= ((((((~(ln_1_nor_33_cse_1 | ln_1_land_17_lpi_1_dfm_1
          | ln_1_land_18_lpi_1_dfm_1 | ln_1_land_19_lpi_1_dfm_1 | ln_1_land_20_lpi_1_dfm_1
          | ln_1_land_21_lpi_1_dfm_1 | ln_1_land_22_lpi_1_dfm_1 | ln_1_land_23_lpi_1_dfm_1
          | ln_1_land_24_lpi_1_dfm_1 | ln_1_land_25_lpi_1_dfm_1 | ln_1_land_26_lpi_1_dfm_1
          | ln_1_land_27_lpi_1_dfm_1 | ln_1_land_28_lpi_1_dfm_1 | ln_1_land_29_lpi_1_dfm_1
          | ln_1_land_30_lpi_1_dfm_1 | ln_1_land_31_lpi_1_dfm_1 | ln_1_land_32_lpi_1_dfm_1
          | ln_1_land_33_lpi_1_dfm_1 | ln_1_land_34_lpi_1_dfm_1 | ln_1_land_35_lpi_1_dfm_1
          | ln_1_land_36_lpi_1_dfm_1 | ln_1_land_37_lpi_1_dfm_1 | ln_1_land_38_lpi_1_dfm_1
          | ln_1_land_39_lpi_1_dfm_1 | ln_1_land_40_lpi_1_dfm_1 | ln_1_land_41_lpi_1_dfm_1
          | ln_1_land_42_lpi_1_dfm_1 | ln_1_land_43_lpi_1_dfm_1 | ln_1_land_44_lpi_1_dfm_1
          | ln_1_land_45_lpi_1_dfm_1 | ln_1_land_46_lpi_1_dfm_1 | ln_1_land_47_lpi_1_dfm_1
          | ln_1_land_48_lpi_1_dfm_1 | ln_1_land_49_lpi_1_dfm_1 | ln_1_if_50_ln_1_if_50_and_seb_1))
          | ln_1_land_51_lpi_1_dfm_1 | ln_1_land_52_lpi_1_dfm_1) & (~(ln_1_land_77_lpi_1_dfm_1
          | ln_1_land_78_lpi_1_dfm_1 | ln_1_land_79_lpi_1_dfm_1 | ln_1_land_80_lpi_1_dfm_1
          | ln_1_land_81_lpi_1_dfm_1 | ln_1_land_82_lpi_1_dfm_1 | ln_1_land_83_lpi_1_dfm_1
          | ln_1_land_84_lpi_1_dfm_1 | ln_1_land_85_lpi_1_dfm_1 | ln_1_land_86_lpi_1_dfm_1
          | ln_1_land_87_lpi_1_dfm_1 | ln_1_land_88_lpi_1_dfm_1 | ln_1_land_89_lpi_1_dfm_1
          | ln_1_land_90_lpi_1_dfm_1 | ln_1_land_91_lpi_1_dfm_1 | ln_1_land_92_lpi_1_dfm_1
          | ln_1_land_93_lpi_1_dfm_1 | ln_1_land_94_lpi_1_dfm_1 | ln_1_land_95_lpi_1_dfm_1
          | ln_1_land_96_lpi_1_dfm_1 | ln_1_land_97_lpi_1_dfm_1 | ln_1_land_114_lpi_1_dfm_1
          | ln_1_land_115_lpi_1_dfm_1 | ln_1_land_116_lpi_1_dfm_1 | ln_1_land_117_lpi_1_dfm_1
          | ln_1_land_118_lpi_1_dfm_1 | ln_1_land_119_lpi_1_dfm_1 | ln_1_land_120_lpi_1_dfm_1
          | ln_1_land_121_lpi_1_dfm_1 | ln_1_land_122_lpi_1_dfm_1 | ln_1_land_123_lpi_1_dfm_1
          | ln_1_land_124_lpi_1_dfm_1 | ln_1_land_125_lpi_1_dfm_1 | ln_1_land_126_lpi_1_dfm_1
          | ln_1_land_127_lpi_1_dfm_1 | ln_1_land_128_lpi_1_dfm_1 | ln_1_land_129_lpi_1_dfm_1
          | ln_1_land_130_lpi_1_dfm_1 | ln_1_land_131_lpi_1_dfm_1 | ln_1_land_132_lpi_1_dfm_1
          | ln_1_land_133_lpi_1_dfm_1 | ln_1_land_134_lpi_1_dfm_1 | ln_1_land_135_lpi_1_dfm_1
          | ln_1_land_136_lpi_1_dfm_1 | ln_1_land_137_lpi_1_dfm_1 | ln_1_land_138_lpi_1_dfm_1
          | ln_1_land_139_lpi_1_dfm_1 | ln_1_land_140_lpi_1_dfm_1))) | ln_1_and_48_ssc_1
          | ln_1_land_54_lpi_1_dfm_1 | ln_1_land_55_lpi_1_dfm_1 | ln_1_land_56_lpi_1_dfm_1
          | ln_1_land_57_lpi_1_dfm_1 | ln_1_land_58_lpi_1_dfm_1 | ln_1_land_59_lpi_1_dfm_1
          | ln_1_land_60_lpi_1_dfm_1 | ln_1_land_61_lpi_1_dfm_1 | ln_1_land_62_lpi_1_dfm_1
          | ln_1_land_63_lpi_1_dfm_1 | ln_1_land_64_lpi_1_dfm_1 | ln_1_land_65_lpi_1_dfm_1
          | ln_1_land_66_lpi_1_dfm_1 | ln_1_land_67_lpi_1_dfm_1 | ln_1_land_68_lpi_1_dfm_1
          | ln_1_land_69_lpi_1_dfm_1 | ln_1_land_70_lpi_1_dfm_1 | ln_1_land_71_lpi_1_dfm_1
          | ln_1_land_72_lpi_1_dfm_1 | ln_1_land_73_lpi_1_dfm_1 | ln_1_land_74_lpi_1_dfm_1
          | ln_1_land_75_lpi_1_dfm_1 | ln_1_land_76_lpi_1_dfm_1 | ln_1_land_98_lpi_1_dfm_1
          | ln_1_land_99_lpi_1_dfm_1 | ln_1_land_100_lpi_1_dfm_1 | ln_1_land_101_lpi_1_dfm_1
          | ln_1_land_102_lpi_1_dfm_1 | ln_1_land_103_lpi_1_dfm_1 | ln_1_land_104_lpi_1_dfm_1
          | ln_1_land_105_lpi_1_dfm_1 | ln_1_land_106_lpi_1_dfm_1 | ln_1_land_107_lpi_1_dfm_1
          | ln_1_land_108_lpi_1_dfm_1 | ln_1_land_109_lpi_1_dfm_1 | ln_1_land_110_lpi_1_dfm_1
          | ln_1_land_111_lpi_1_dfm_1 | ln_1_land_112_lpi_1_dfm_1 | ln_1_land_113_lpi_1_dfm_1
          | ln_1_land_141_lpi_1_dfm_1 | ln_1_land_142_lpi_1_dfm_1 | ln_1_and_138_ssc_1
          | ln_1_land_144_lpi_1_dfm_1) & (~(ln_1_land_172_lpi_1_dfm_1 | ln_1_land_173_lpi_1_dfm_1
          | ln_1_land_174_lpi_1_dfm_1 | ln_1_land_175_lpi_1_dfm_1 | ln_1_land_176_lpi_1_dfm_1
          | ln_1_land_177_lpi_1_dfm_1 | ln_1_land_178_lpi_1_dfm_1 | ln_1_land_179_lpi_1_dfm_1
          | ln_1_land_180_lpi_1_dfm_1 | ln_1_land_181_lpi_1_dfm_1 | ln_1_land_182_lpi_1_dfm_1
          | ln_1_land_183_lpi_1_dfm_1 | ln_1_land_184_lpi_1_dfm_1 | ln_1_land_185_lpi_1_dfm_1
          | ln_1_land_186_lpi_1_dfm_1 | ln_1_land_187_lpi_1_dfm_1 | ln_1_land_188_lpi_1_dfm_1
          | ln_1_land_189_lpi_1_dfm_1 | ln_1_land_190_lpi_1_dfm_1 | ln_1_land_191_lpi_1_dfm_1
          | ln_1_land_192_lpi_1_dfm_1 | ln_1_land_193_lpi_1_dfm_1 | ln_1_land_194_lpi_1_dfm_1
          | ln_1_land_214_lpi_1_dfm_1 | ln_1_land_215_lpi_1_dfm_1 | ln_1_land_216_lpi_1_dfm_1
          | ln_1_land_217_lpi_1_dfm_1 | ln_1_land_218_lpi_1_dfm_1 | ln_1_land_219_lpi_1_dfm_1
          | ln_1_land_220_lpi_1_dfm_1 | ln_1_land_221_lpi_1_dfm_1 | ln_1_land_222_lpi_1_dfm_1
          | ln_1_land_223_lpi_1_dfm_1 | ln_1_land_224_lpi_1_dfm_1 | ln_1_land_225_lpi_1_dfm_1
          | ln_1_land_226_lpi_1_dfm_1 | ln_1_land_227_lpi_1_dfm_1 | ln_1_land_228_lpi_1_dfm_1
          | ln_1_land_240_lpi_1_dfm_1 | ln_1_land_241_lpi_1_dfm_1 | ln_1_land_242_lpi_1_dfm_1
          | ln_1_land_243_lpi_1_dfm_1 | ln_1_land_244_lpi_1_dfm_1))) | ln_1_and_140_ssc_1
          | ln_1_land_146_lpi_1_dfm_1 | ln_1_land_147_lpi_1_dfm_1 | ln_1_land_148_lpi_1_dfm_1
          | ln_1_land_149_lpi_1_dfm_1 | ln_1_land_150_lpi_1_dfm_1 | ln_1_land_151_lpi_1_dfm_1
          | ln_1_land_152_lpi_1_dfm_1 | ln_1_land_153_lpi_1_dfm_1 | ln_1_land_154_lpi_1_dfm_1
          | ln_1_land_155_lpi_1_dfm_1 | ln_1_land_156_lpi_1_dfm_1 | ln_1_land_157_lpi_1_dfm_1
          | ln_1_land_158_lpi_1_dfm_1 | ln_1_land_159_lpi_1_dfm_1 | ln_1_land_160_lpi_1_dfm_1
          | ln_1_land_161_lpi_1_dfm_1 | ln_1_land_162_lpi_1_dfm_1 | ln_1_land_163_lpi_1_dfm_1
          | ln_1_land_164_lpi_1_dfm_1 | ln_1_land_165_lpi_1_dfm_1 | ln_1_land_166_lpi_1_dfm_1
          | ln_1_land_167_lpi_1_dfm_1 | ln_1_land_168_lpi_1_dfm_1 | ln_1_land_169_lpi_1_dfm_1
          | ln_1_land_170_lpi_1_dfm_1 | ln_1_land_171_lpi_1_dfm_1 | ln_1_land_195_lpi_1_dfm_1
          | ln_1_land_196_lpi_1_dfm_1 | ln_1_land_197_lpi_1_dfm_1 | ln_1_land_198_lpi_1_dfm_1
          | ln_1_land_199_lpi_1_dfm_1 | ln_1_land_200_lpi_1_dfm_1 | ln_1_land_201_lpi_1_dfm_1
          | ln_1_land_202_lpi_1_dfm_1 | ln_1_land_203_lpi_1_dfm_1 | ln_1_land_204_lpi_1_dfm_1
          | ln_1_land_205_lpi_1_dfm_1 | ln_1_land_206_lpi_1_dfm_1 | ln_1_land_207_lpi_1_dfm_1
          | ln_1_land_208_lpi_1_dfm_1 | ln_1_land_209_lpi_1_dfm_1 | ln_1_land_210_lpi_1_dfm_1
          | ln_1_land_211_lpi_1_dfm_1 | ln_1_land_212_lpi_1_dfm_1 | ln_1_land_213_lpi_1_dfm_1
          | ln_1_land_229_lpi_1_dfm_1 | ln_1_land_230_lpi_1_dfm_1 | ln_1_land_231_lpi_1_dfm_1
          | ln_1_land_232_lpi_1_dfm_1 | ln_1_land_233_lpi_1_dfm_1 | ln_1_land_234_lpi_1_dfm_1
          | ln_1_land_235_lpi_1_dfm_1 | ln_1_land_236_lpi_1_dfm_1 | ln_1_land_237_lpi_1_dfm_1
          | ln_1_land_238_lpi_1_dfm_1 | ln_1_land_239_lpi_1_dfm_1) & (~(ln_1_and_240_ssc_1_1
          | ln_1_land_246_lpi_1_dfm_1 | ln_1_land_247_lpi_1_dfm_1 | ln_1_land_249_lpi_1_dfm_1
          | ln_1_land_250_lpi_1_dfm_1 | ln_1_land_252_lpi_1_dfm_1_1));
      ln_1_ln_1_mux1h_118_psp_1_8 <= (((((~(((~((~(ln_1_nor_5_cse_1 | ln_1_and_2_ssc_1))
          | ln_1_land_6_lpi_1_dfm_1)) & (~(ln_1_land_17_lpi_1_dfm_1 | ln_1_land_18_lpi_1_dfm_1
          | ln_1_land_19_lpi_1_dfm_1 | ln_1_land_20_lpi_1_dfm_1 | ln_1_land_21_lpi_1_dfm_1
          | ln_1_land_22_lpi_1_dfm_1 | ln_1_land_23_lpi_1_dfm_1 | ln_1_land_24_lpi_1_dfm_1
          | ln_1_land_25_lpi_1_dfm_1 | ln_1_land_26_lpi_1_dfm_1 | ln_1_land_27_lpi_1_dfm_1
          | ln_1_land_28_lpi_1_dfm_1 | ln_1_land_29_lpi_1_dfm_1 | ln_1_land_30_lpi_1_dfm_1
          | ln_1_land_31_lpi_1_dfm_1 | ln_1_land_32_lpi_1_dfm_1 | ln_1_land_33_lpi_1_dfm_1
          | ln_1_land_34_lpi_1_dfm_1))) | ln_1_and_4_ssc_1 | ln_1_land_8_lpi_1_dfm_1
          | ln_1_land_9_lpi_1_dfm_1 | ln_1_land_10_lpi_1_dfm_1 | ln_1_land_11_lpi_1_dfm_1
          | ln_1_land_12_lpi_1_dfm_1 | ln_1_land_13_lpi_1_dfm_1 | ln_1_land_14_lpi_1_dfm_1
          | ln_1_land_15_lpi_1_dfm_1 | ln_1_land_16_lpi_1_dfm_1 | ln_1_land_35_lpi_1_dfm_1
          | ln_1_land_36_lpi_1_dfm_1 | ln_1_land_37_lpi_1_dfm_1 | ln_1_land_38_lpi_1_dfm_1
          | ln_1_land_39_lpi_1_dfm_1 | ln_1_land_40_lpi_1_dfm_1 | ln_1_land_41_lpi_1_dfm_1
          | ln_1_land_42_lpi_1_dfm_1 | ln_1_land_43_lpi_1_dfm_1 | ln_1_land_44_lpi_1_dfm_1
          | ln_1_land_45_lpi_1_dfm_1 | ln_1_land_46_lpi_1_dfm_1 | ln_1_land_47_lpi_1_dfm_1
          | ln_1_land_48_lpi_1_dfm_1 | ln_1_land_49_lpi_1_dfm_1 | ln_1_if_50_ln_1_if_50_and_seb_1))
          | ln_1_land_51_lpi_1_dfm_1 | ln_1_land_52_lpi_1_dfm_1) & (~(ln_1_land_65_lpi_1_dfm_1
          | ln_1_land_66_lpi_1_dfm_1 | ln_1_land_67_lpi_1_dfm_1 | ln_1_land_68_lpi_1_dfm_1
          | ln_1_land_69_lpi_1_dfm_1 | ln_1_land_70_lpi_1_dfm_1 | ln_1_land_71_lpi_1_dfm_1
          | ln_1_land_72_lpi_1_dfm_1 | ln_1_land_73_lpi_1_dfm_1 | ln_1_land_74_lpi_1_dfm_1
          | ln_1_land_75_lpi_1_dfm_1 | ln_1_land_76_lpi_1_dfm_1 | ln_1_land_88_lpi_1_dfm_1
          | ln_1_land_89_lpi_1_dfm_1 | ln_1_land_90_lpi_1_dfm_1 | ln_1_land_91_lpi_1_dfm_1
          | ln_1_land_92_lpi_1_dfm_1 | ln_1_land_93_lpi_1_dfm_1 | ln_1_land_94_lpi_1_dfm_1
          | ln_1_land_95_lpi_1_dfm_1 | ln_1_land_96_lpi_1_dfm_1 | ln_1_land_97_lpi_1_dfm_1
          | ln_1_land_106_lpi_1_dfm_1 | ln_1_land_107_lpi_1_dfm_1 | ln_1_land_108_lpi_1_dfm_1
          | ln_1_land_109_lpi_1_dfm_1 | ln_1_land_110_lpi_1_dfm_1 | ln_1_land_111_lpi_1_dfm_1
          | ln_1_land_112_lpi_1_dfm_1 | ln_1_land_113_lpi_1_dfm_1 | ln_1_land_122_lpi_1_dfm_1
          | ln_1_land_123_lpi_1_dfm_1 | ln_1_land_124_lpi_1_dfm_1 | ln_1_land_125_lpi_1_dfm_1
          | ln_1_land_126_lpi_1_dfm_1 | ln_1_land_127_lpi_1_dfm_1 | ln_1_land_128_lpi_1_dfm_1
          | ln_1_land_129_lpi_1_dfm_1 | ln_1_land_130_lpi_1_dfm_1 | ln_1_land_131_lpi_1_dfm_1
          | ln_1_land_132_lpi_1_dfm_1 | ln_1_land_133_lpi_1_dfm_1 | ln_1_land_134_lpi_1_dfm_1
          | ln_1_land_135_lpi_1_dfm_1 | ln_1_land_136_lpi_1_dfm_1 | ln_1_land_137_lpi_1_dfm_1
          | ln_1_land_138_lpi_1_dfm_1 | ln_1_land_139_lpi_1_dfm_1 | ln_1_land_140_lpi_1_dfm_1)))
          | ln_1_and_48_ssc_1 | ln_1_land_54_lpi_1_dfm_1 | ln_1_land_55_lpi_1_dfm_1
          | ln_1_land_56_lpi_1_dfm_1 | ln_1_land_57_lpi_1_dfm_1 | ln_1_land_58_lpi_1_dfm_1
          | ln_1_land_59_lpi_1_dfm_1 | ln_1_land_60_lpi_1_dfm_1 | ln_1_land_61_lpi_1_dfm_1
          | ln_1_land_62_lpi_1_dfm_1 | ln_1_land_63_lpi_1_dfm_1 | ln_1_land_64_lpi_1_dfm_1
          | ln_1_land_77_lpi_1_dfm_1 | ln_1_land_78_lpi_1_dfm_1 | ln_1_land_79_lpi_1_dfm_1
          | ln_1_land_80_lpi_1_dfm_1 | ln_1_land_81_lpi_1_dfm_1 | ln_1_land_82_lpi_1_dfm_1
          | ln_1_land_83_lpi_1_dfm_1 | ln_1_land_84_lpi_1_dfm_1 | ln_1_land_85_lpi_1_dfm_1
          | ln_1_land_86_lpi_1_dfm_1 | ln_1_land_87_lpi_1_dfm_1 | ln_1_land_98_lpi_1_dfm_1
          | ln_1_land_99_lpi_1_dfm_1 | ln_1_land_100_lpi_1_dfm_1 | ln_1_land_101_lpi_1_dfm_1
          | ln_1_land_102_lpi_1_dfm_1 | ln_1_land_103_lpi_1_dfm_1 | ln_1_land_104_lpi_1_dfm_1
          | ln_1_land_105_lpi_1_dfm_1 | ln_1_land_114_lpi_1_dfm_1 | ln_1_land_115_lpi_1_dfm_1
          | ln_1_land_116_lpi_1_dfm_1 | ln_1_land_117_lpi_1_dfm_1 | ln_1_land_118_lpi_1_dfm_1
          | ln_1_land_119_lpi_1_dfm_1 | ln_1_land_120_lpi_1_dfm_1 | ln_1_land_121_lpi_1_dfm_1
          | ln_1_land_141_lpi_1_dfm_1 | ln_1_land_142_lpi_1_dfm_1 | ln_1_and_138_ssc_1
          | ln_1_land_144_lpi_1_dfm_1) & (~(ln_1_land_157_lpi_1_dfm_1 | ln_1_land_158_lpi_1_dfm_1
          | ln_1_land_159_lpi_1_dfm_1 | ln_1_land_160_lpi_1_dfm_1 | ln_1_land_161_lpi_1_dfm_1
          | ln_1_land_162_lpi_1_dfm_1 | ln_1_land_163_lpi_1_dfm_1 | ln_1_land_164_lpi_1_dfm_1
          | ln_1_land_165_lpi_1_dfm_1 | ln_1_land_166_lpi_1_dfm_1 | ln_1_land_167_lpi_1_dfm_1
          | ln_1_land_168_lpi_1_dfm_1 | ln_1_land_169_lpi_1_dfm_1 | ln_1_land_170_lpi_1_dfm_1
          | ln_1_land_171_lpi_1_dfm_1 | ln_1_land_184_lpi_1_dfm_1 | ln_1_land_185_lpi_1_dfm_1
          | ln_1_land_186_lpi_1_dfm_1 | ln_1_land_187_lpi_1_dfm_1 | ln_1_land_188_lpi_1_dfm_1
          | ln_1_land_189_lpi_1_dfm_1 | ln_1_land_190_lpi_1_dfm_1 | ln_1_land_191_lpi_1_dfm_1
          | ln_1_land_192_lpi_1_dfm_1 | ln_1_land_193_lpi_1_dfm_1 | ln_1_land_194_lpi_1_dfm_1
          | ln_1_land_205_lpi_1_dfm_1 | ln_1_land_206_lpi_1_dfm_1 | ln_1_land_207_lpi_1_dfm_1
          | ln_1_land_208_lpi_1_dfm_1 | ln_1_land_209_lpi_1_dfm_1 | ln_1_land_210_lpi_1_dfm_1
          | ln_1_land_211_lpi_1_dfm_1 | ln_1_land_212_lpi_1_dfm_1 | ln_1_land_213_lpi_1_dfm_1
          | ln_1_land_222_lpi_1_dfm_1 | ln_1_land_223_lpi_1_dfm_1 | ln_1_land_224_lpi_1_dfm_1
          | ln_1_land_225_lpi_1_dfm_1 | ln_1_land_226_lpi_1_dfm_1 | ln_1_land_227_lpi_1_dfm_1
          | ln_1_land_228_lpi_1_dfm_1 | ln_1_land_235_lpi_1_dfm_1 | ln_1_land_236_lpi_1_dfm_1
          | ln_1_land_237_lpi_1_dfm_1 | ln_1_land_238_lpi_1_dfm_1 | ln_1_land_239_lpi_1_dfm_1
          | ln_1_land_244_lpi_1_dfm_1))) | ln_1_and_140_ssc_1 | ln_1_land_146_lpi_1_dfm_1
          | ln_1_land_147_lpi_1_dfm_1 | ln_1_land_148_lpi_1_dfm_1 | ln_1_land_149_lpi_1_dfm_1
          | ln_1_land_150_lpi_1_dfm_1 | ln_1_land_151_lpi_1_dfm_1 | ln_1_land_152_lpi_1_dfm_1
          | ln_1_land_153_lpi_1_dfm_1 | ln_1_land_154_lpi_1_dfm_1 | ln_1_land_155_lpi_1_dfm_1
          | ln_1_land_156_lpi_1_dfm_1 | ln_1_land_172_lpi_1_dfm_1 | ln_1_land_173_lpi_1_dfm_1
          | ln_1_land_174_lpi_1_dfm_1 | ln_1_land_175_lpi_1_dfm_1 | ln_1_land_176_lpi_1_dfm_1
          | ln_1_land_177_lpi_1_dfm_1 | ln_1_land_178_lpi_1_dfm_1 | ln_1_land_179_lpi_1_dfm_1
          | ln_1_land_180_lpi_1_dfm_1 | ln_1_land_181_lpi_1_dfm_1 | ln_1_land_182_lpi_1_dfm_1
          | ln_1_land_183_lpi_1_dfm_1 | ln_1_land_195_lpi_1_dfm_1 | ln_1_land_196_lpi_1_dfm_1
          | ln_1_land_197_lpi_1_dfm_1 | ln_1_land_198_lpi_1_dfm_1 | ln_1_land_199_lpi_1_dfm_1
          | ln_1_land_200_lpi_1_dfm_1 | ln_1_land_201_lpi_1_dfm_1 | ln_1_land_202_lpi_1_dfm_1
          | ln_1_land_203_lpi_1_dfm_1 | ln_1_land_204_lpi_1_dfm_1 | ln_1_land_214_lpi_1_dfm_1
          | ln_1_land_215_lpi_1_dfm_1 | ln_1_land_216_lpi_1_dfm_1 | ln_1_land_217_lpi_1_dfm_1
          | ln_1_land_218_lpi_1_dfm_1 | ln_1_land_219_lpi_1_dfm_1 | ln_1_land_220_lpi_1_dfm_1
          | ln_1_land_221_lpi_1_dfm_1 | ln_1_land_229_lpi_1_dfm_1 | ln_1_land_230_lpi_1_dfm_1
          | ln_1_land_231_lpi_1_dfm_1 | ln_1_land_232_lpi_1_dfm_1 | ln_1_land_233_lpi_1_dfm_1
          | ln_1_land_234_lpi_1_dfm_1 | ln_1_land_240_lpi_1_dfm_1 | ln_1_land_241_lpi_1_dfm_1
          | ln_1_land_242_lpi_1_dfm_1 | ln_1_land_243_lpi_1_dfm_1;
      ln_1_ln_1_mux1h_118_psp_1_7 <= (((((~(((~(ln_1_ln_1_ln_1_nor_8_cse_1 & ln_1_nor_1_cse_1))
          & (~(ln_1_land_17_lpi_1_dfm_1 | ln_1_land_18_lpi_1_dfm_1 | ln_1_land_19_lpi_1_dfm_1
          | ln_1_land_20_lpi_1_dfm_1 | ln_1_land_21_lpi_1_dfm_1 | ln_1_land_22_lpi_1_dfm_1
          | ln_1_land_23_lpi_1_dfm_1 | ln_1_land_24_lpi_1_dfm_1 | ln_1_land_25_lpi_1_dfm_1
          | ln_1_land_35_lpi_1_dfm_1 | ln_1_land_36_lpi_1_dfm_1 | ln_1_land_37_lpi_1_dfm_1
          | ln_1_land_38_lpi_1_dfm_1 | ln_1_land_39_lpi_1_dfm_1 | ln_1_land_40_lpi_1_dfm_1
          | ln_1_land_41_lpi_1_dfm_1 | ln_1_land_42_lpi_1_dfm_1))) | ln_1_and_4_ssc_1
          | ln_1_land_8_lpi_1_dfm_1 | ln_1_land_9_lpi_1_dfm_1 | ln_1_land_10_lpi_1_dfm_1
          | ln_1_land_11_lpi_1_dfm_1 | ln_1_land_12_lpi_1_dfm_1 | ln_1_land_13_lpi_1_dfm_1
          | ln_1_land_14_lpi_1_dfm_1 | ln_1_land_15_lpi_1_dfm_1 | ln_1_land_16_lpi_1_dfm_1
          | ln_1_land_26_lpi_1_dfm_1 | ln_1_land_27_lpi_1_dfm_1 | ln_1_land_28_lpi_1_dfm_1
          | ln_1_land_29_lpi_1_dfm_1 | ln_1_land_30_lpi_1_dfm_1 | ln_1_land_31_lpi_1_dfm_1
          | ln_1_land_32_lpi_1_dfm_1 | ln_1_land_33_lpi_1_dfm_1 | ln_1_land_34_lpi_1_dfm_1
          | ln_1_land_43_lpi_1_dfm_1 | ln_1_land_44_lpi_1_dfm_1 | ln_1_land_45_lpi_1_dfm_1
          | ln_1_land_46_lpi_1_dfm_1 | ln_1_land_47_lpi_1_dfm_1 | ln_1_land_48_lpi_1_dfm_1
          | ln_1_land_49_lpi_1_dfm_1 | ln_1_if_50_ln_1_if_50_and_seb_1)) | ln_1_land_51_lpi_1_dfm_1
          | ln_1_land_52_lpi_1_dfm_1) & (~(ln_1_land_58_lpi_1_dfm_1 | ln_1_land_59_lpi_1_dfm_1
          | ln_1_land_60_lpi_1_dfm_1 | ln_1_land_61_lpi_1_dfm_1 | ln_1_land_62_lpi_1_dfm_1
          | ln_1_land_63_lpi_1_dfm_1 | ln_1_land_64_lpi_1_dfm_1 | ln_1_land_71_lpi_1_dfm_1
          | ln_1_land_72_lpi_1_dfm_1 | ln_1_land_73_lpi_1_dfm_1 | ln_1_land_74_lpi_1_dfm_1
          | ln_1_land_75_lpi_1_dfm_1 | ln_1_land_76_lpi_1_dfm_1 | ln_1_land_83_lpi_1_dfm_1
          | ln_1_land_84_lpi_1_dfm_1 | ln_1_land_85_lpi_1_dfm_1 | ln_1_land_86_lpi_1_dfm_1
          | ln_1_land_87_lpi_1_dfm_1 | ln_1_land_93_lpi_1_dfm_1 | ln_1_land_94_lpi_1_dfm_1
          | ln_1_land_95_lpi_1_dfm_1 | ln_1_land_96_lpi_1_dfm_1 | ln_1_land_97_lpi_1_dfm_1
          | ln_1_land_102_lpi_1_dfm_1 | ln_1_land_103_lpi_1_dfm_1 | ln_1_land_104_lpi_1_dfm_1
          | ln_1_land_105_lpi_1_dfm_1 | ln_1_land_110_lpi_1_dfm_1 | ln_1_land_111_lpi_1_dfm_1
          | ln_1_land_112_lpi_1_dfm_1 | ln_1_land_113_lpi_1_dfm_1 | ln_1_land_117_lpi_1_dfm_1
          | ln_1_land_118_lpi_1_dfm_1 | ln_1_land_119_lpi_1_dfm_1 | ln_1_land_120_lpi_1_dfm_1
          | ln_1_land_121_lpi_1_dfm_1 | ln_1_land_132_lpi_1_dfm_1 | ln_1_land_133_lpi_1_dfm_1
          | ln_1_land_134_lpi_1_dfm_1 | ln_1_land_135_lpi_1_dfm_1 | ln_1_land_136_lpi_1_dfm_1
          | ln_1_land_137_lpi_1_dfm_1 | ln_1_land_138_lpi_1_dfm_1 | ln_1_land_139_lpi_1_dfm_1
          | ln_1_land_140_lpi_1_dfm_1))) | ln_1_and_48_ssc_1 | ln_1_land_54_lpi_1_dfm_1
          | ln_1_land_55_lpi_1_dfm_1 | ln_1_land_56_lpi_1_dfm_1 | ln_1_land_57_lpi_1_dfm_1
          | ln_1_land_65_lpi_1_dfm_1 | ln_1_land_66_lpi_1_dfm_1 | ln_1_land_67_lpi_1_dfm_1
          | ln_1_land_68_lpi_1_dfm_1 | ln_1_land_69_lpi_1_dfm_1 | ln_1_land_70_lpi_1_dfm_1
          | ln_1_land_77_lpi_1_dfm_1 | ln_1_land_78_lpi_1_dfm_1 | ln_1_land_79_lpi_1_dfm_1
          | ln_1_land_80_lpi_1_dfm_1 | ln_1_land_81_lpi_1_dfm_1 | ln_1_land_82_lpi_1_dfm_1
          | ln_1_land_88_lpi_1_dfm_1 | ln_1_land_89_lpi_1_dfm_1 | ln_1_land_90_lpi_1_dfm_1
          | ln_1_land_91_lpi_1_dfm_1 | ln_1_land_92_lpi_1_dfm_1 | ln_1_land_98_lpi_1_dfm_1
          | ln_1_land_99_lpi_1_dfm_1 | ln_1_land_100_lpi_1_dfm_1 | ln_1_land_101_lpi_1_dfm_1
          | ln_1_land_106_lpi_1_dfm_1 | ln_1_land_107_lpi_1_dfm_1 | ln_1_land_108_lpi_1_dfm_1
          | ln_1_land_109_lpi_1_dfm_1 | ln_1_land_114_lpi_1_dfm_1 | ln_1_land_115_lpi_1_dfm_1
          | ln_1_land_116_lpi_1_dfm_1 | ln_1_land_122_lpi_1_dfm_1 | ln_1_land_123_lpi_1_dfm_1
          | ln_1_land_124_lpi_1_dfm_1 | ln_1_land_125_lpi_1_dfm_1 | ln_1_land_126_lpi_1_dfm_1
          | ln_1_land_127_lpi_1_dfm_1 | ln_1_land_128_lpi_1_dfm_1 | ln_1_land_129_lpi_1_dfm_1
          | ln_1_land_130_lpi_1_dfm_1 | ln_1_land_131_lpi_1_dfm_1 | ln_1_land_141_lpi_1_dfm_1
          | ln_1_land_142_lpi_1_dfm_1 | ln_1_and_138_ssc_1 | ln_1_land_144_lpi_1_dfm_1)
          & (~(ln_1_land_149_lpi_1_dfm_1 | ln_1_land_150_lpi_1_dfm_1 | ln_1_land_151_lpi_1_dfm_1
          | ln_1_land_152_lpi_1_dfm_1 | ln_1_land_153_lpi_1_dfm_1 | ln_1_land_154_lpi_1_dfm_1
          | ln_1_land_155_lpi_1_dfm_1 | ln_1_land_156_lpi_1_dfm_1 | ln_1_land_165_lpi_1_dfm_1
          | ln_1_land_166_lpi_1_dfm_1 | ln_1_land_167_lpi_1_dfm_1 | ln_1_land_168_lpi_1_dfm_1
          | ln_1_land_169_lpi_1_dfm_1 | ln_1_land_170_lpi_1_dfm_1 | ln_1_land_171_lpi_1_dfm_1
          | ln_1_land_178_lpi_1_dfm_1 | ln_1_land_179_lpi_1_dfm_1 | ln_1_land_180_lpi_1_dfm_1
          | ln_1_land_181_lpi_1_dfm_1 | ln_1_land_182_lpi_1_dfm_1 | ln_1_land_183_lpi_1_dfm_1
          | ln_1_land_190_lpi_1_dfm_1 | ln_1_land_191_lpi_1_dfm_1 | ln_1_land_192_lpi_1_dfm_1
          | ln_1_land_193_lpi_1_dfm_1 | ln_1_land_194_lpi_1_dfm_1 | ln_1_land_201_lpi_1_dfm_1
          | ln_1_land_202_lpi_1_dfm_1 | ln_1_land_203_lpi_1_dfm_1 | ln_1_land_204_lpi_1_dfm_1
          | ln_1_land_210_lpi_1_dfm_1 | ln_1_land_211_lpi_1_dfm_1 | ln_1_land_212_lpi_1_dfm_1
          | ln_1_land_213_lpi_1_dfm_1 | ln_1_land_218_lpi_1_dfm_1 | ln_1_land_219_lpi_1_dfm_1
          | ln_1_land_220_lpi_1_dfm_1 | ln_1_land_221_lpi_1_dfm_1 | ln_1_land_225_lpi_1_dfm_1
          | ln_1_land_226_lpi_1_dfm_1 | ln_1_land_227_lpi_1_dfm_1 | ln_1_land_228_lpi_1_dfm_1
          | ln_1_land_232_lpi_1_dfm_1 | ln_1_land_233_lpi_1_dfm_1 | ln_1_land_234_lpi_1_dfm_1
          | ln_1_land_237_lpi_1_dfm_1 | ln_1_land_238_lpi_1_dfm_1 | ln_1_land_239_lpi_1_dfm_1
          | ln_1_land_242_lpi_1_dfm_1 | ln_1_land_243_lpi_1_dfm_1))) | ln_1_and_140_ssc_1
          | ln_1_land_146_lpi_1_dfm_1 | ln_1_land_147_lpi_1_dfm_1 | ln_1_land_148_lpi_1_dfm_1
          | ln_1_land_157_lpi_1_dfm_1 | ln_1_land_158_lpi_1_dfm_1 | ln_1_land_159_lpi_1_dfm_1
          | ln_1_land_160_lpi_1_dfm_1 | ln_1_land_161_lpi_1_dfm_1 | ln_1_land_162_lpi_1_dfm_1
          | ln_1_land_163_lpi_1_dfm_1 | ln_1_land_164_lpi_1_dfm_1 | ln_1_land_172_lpi_1_dfm_1
          | ln_1_land_173_lpi_1_dfm_1 | ln_1_land_174_lpi_1_dfm_1 | ln_1_land_175_lpi_1_dfm_1
          | ln_1_land_176_lpi_1_dfm_1 | ln_1_land_177_lpi_1_dfm_1 | ln_1_land_184_lpi_1_dfm_1
          | ln_1_land_185_lpi_1_dfm_1 | ln_1_land_186_lpi_1_dfm_1 | ln_1_land_187_lpi_1_dfm_1
          | ln_1_land_188_lpi_1_dfm_1 | ln_1_land_189_lpi_1_dfm_1 | ln_1_land_195_lpi_1_dfm_1
          | ln_1_land_196_lpi_1_dfm_1 | ln_1_land_197_lpi_1_dfm_1 | ln_1_land_198_lpi_1_dfm_1
          | ln_1_land_199_lpi_1_dfm_1 | ln_1_land_200_lpi_1_dfm_1 | ln_1_land_205_lpi_1_dfm_1
          | ln_1_land_206_lpi_1_dfm_1 | ln_1_land_207_lpi_1_dfm_1 | ln_1_land_208_lpi_1_dfm_1
          | ln_1_land_209_lpi_1_dfm_1 | ln_1_land_214_lpi_1_dfm_1 | ln_1_land_215_lpi_1_dfm_1
          | ln_1_land_216_lpi_1_dfm_1 | ln_1_land_217_lpi_1_dfm_1 | ln_1_land_222_lpi_1_dfm_1
          | ln_1_land_223_lpi_1_dfm_1 | ln_1_land_224_lpi_1_dfm_1 | ln_1_land_229_lpi_1_dfm_1
          | ln_1_land_230_lpi_1_dfm_1 | ln_1_land_231_lpi_1_dfm_1 | ln_1_land_235_lpi_1_dfm_1
          | ln_1_land_236_lpi_1_dfm_1 | ln_1_land_240_lpi_1_dfm_1 | ln_1_land_241_lpi_1_dfm_1
          | ln_1_land_244_lpi_1_dfm_1;
      ln_1_ln_1_mux1h_118_psp_1_6 <= (((((~(ln_1_nor_33_cse_1 | ln_1_land_12_lpi_1_dfm_1
          | ln_1_land_13_lpi_1_dfm_1 | ln_1_land_14_lpi_1_dfm_1 | ln_1_land_15_lpi_1_dfm_1
          | ln_1_land_16_lpi_1_dfm_1 | ln_1_land_21_lpi_1_dfm_1 | ln_1_land_22_lpi_1_dfm_1
          | ln_1_land_23_lpi_1_dfm_1 | ln_1_land_24_lpi_1_dfm_1 | ln_1_land_25_lpi_1_dfm_1
          | ln_1_land_30_lpi_1_dfm_1 | ln_1_land_31_lpi_1_dfm_1 | ln_1_land_32_lpi_1_dfm_1
          | ln_1_land_33_lpi_1_dfm_1 | ln_1_land_34_lpi_1_dfm_1 | ln_1_land_39_lpi_1_dfm_1
          | ln_1_land_40_lpi_1_dfm_1 | ln_1_land_41_lpi_1_dfm_1 | ln_1_land_42_lpi_1_dfm_1
          | ln_1_land_47_lpi_1_dfm_1 | ln_1_land_48_lpi_1_dfm_1 | ln_1_land_49_lpi_1_dfm_1
          | ln_1_if_50_ln_1_if_50_and_seb_1)) | ln_1_land_51_lpi_1_dfm_1 | ln_1_land_52_lpi_1_dfm_1)
          & (~(ln_1_land_54_lpi_1_dfm_1 | ln_1_land_55_lpi_1_dfm_1 | ln_1_land_56_lpi_1_dfm_1
          | ln_1_land_57_lpi_1_dfm_1 | ln_1_land_61_lpi_1_dfm_1 | ln_1_land_62_lpi_1_dfm_1
          | ln_1_land_63_lpi_1_dfm_1 | ln_1_land_64_lpi_1_dfm_1 | ln_1_land_68_lpi_1_dfm_1
          | ln_1_land_69_lpi_1_dfm_1 | ln_1_land_70_lpi_1_dfm_1 | ln_1_land_74_lpi_1_dfm_1
          | ln_1_land_75_lpi_1_dfm_1 | ln_1_land_76_lpi_1_dfm_1 | ln_1_land_80_lpi_1_dfm_1
          | ln_1_land_81_lpi_1_dfm_1 | ln_1_land_82_lpi_1_dfm_1 | ln_1_land_85_lpi_1_dfm_1
          | ln_1_land_86_lpi_1_dfm_1 | ln_1_land_87_lpi_1_dfm_1 | ln_1_land_91_lpi_1_dfm_1
          | ln_1_land_92_lpi_1_dfm_1 | ln_1_land_95_lpi_1_dfm_1 | ln_1_land_96_lpi_1_dfm_1
          | ln_1_land_97_lpi_1_dfm_1 | ln_1_land_100_lpi_1_dfm_1 | ln_1_land_101_lpi_1_dfm_1
          | ln_1_land_104_lpi_1_dfm_1 | ln_1_land_105_lpi_1_dfm_1 | ln_1_land_108_lpi_1_dfm_1
          | ln_1_land_109_lpi_1_dfm_1 | ln_1_land_112_lpi_1_dfm_1 | ln_1_land_113_lpi_1_dfm_1
          | ln_1_land_116_lpi_1_dfm_1 | ln_1_land_119_lpi_1_dfm_1 | ln_1_land_120_lpi_1_dfm_1
          | ln_1_land_121_lpi_1_dfm_1 | ln_1_land_127_lpi_1_dfm_1 | ln_1_land_128_lpi_1_dfm_1
          | ln_1_land_129_lpi_1_dfm_1 | ln_1_land_130_lpi_1_dfm_1 | ln_1_land_131_lpi_1_dfm_1
          | ln_1_land_137_lpi_1_dfm_1 | ln_1_land_138_lpi_1_dfm_1 | ln_1_land_139_lpi_1_dfm_1
          | ln_1_land_140_lpi_1_dfm_1))) | ln_1_and_48_ssc_1 | ln_1_land_58_lpi_1_dfm_1
          | ln_1_land_59_lpi_1_dfm_1 | ln_1_land_60_lpi_1_dfm_1 | ln_1_land_65_lpi_1_dfm_1
          | ln_1_land_66_lpi_1_dfm_1 | ln_1_land_67_lpi_1_dfm_1 | ln_1_land_71_lpi_1_dfm_1
          | ln_1_land_72_lpi_1_dfm_1 | ln_1_land_73_lpi_1_dfm_1 | ln_1_land_77_lpi_1_dfm_1
          | ln_1_land_78_lpi_1_dfm_1 | ln_1_land_79_lpi_1_dfm_1 | ln_1_land_83_lpi_1_dfm_1
          | ln_1_land_84_lpi_1_dfm_1 | ln_1_land_88_lpi_1_dfm_1 | ln_1_land_89_lpi_1_dfm_1
          | ln_1_land_90_lpi_1_dfm_1 | ln_1_land_93_lpi_1_dfm_1 | ln_1_land_94_lpi_1_dfm_1
          | ln_1_land_98_lpi_1_dfm_1 | ln_1_land_99_lpi_1_dfm_1 | ln_1_land_102_lpi_1_dfm_1
          | ln_1_land_103_lpi_1_dfm_1 | ln_1_land_106_lpi_1_dfm_1 | ln_1_land_107_lpi_1_dfm_1
          | ln_1_land_110_lpi_1_dfm_1 | ln_1_land_111_lpi_1_dfm_1 | ln_1_land_114_lpi_1_dfm_1
          | ln_1_land_115_lpi_1_dfm_1 | ln_1_land_117_lpi_1_dfm_1 | ln_1_land_118_lpi_1_dfm_1
          | ln_1_land_122_lpi_1_dfm_1 | ln_1_land_123_lpi_1_dfm_1 | ln_1_land_124_lpi_1_dfm_1
          | ln_1_land_125_lpi_1_dfm_1 | ln_1_land_126_lpi_1_dfm_1 | ln_1_land_132_lpi_1_dfm_1
          | ln_1_land_133_lpi_1_dfm_1 | ln_1_land_134_lpi_1_dfm_1 | ln_1_land_135_lpi_1_dfm_1
          | ln_1_land_136_lpi_1_dfm_1 | ln_1_land_141_lpi_1_dfm_1 | ln_1_land_142_lpi_1_dfm_1
          | ln_1_and_138_ssc_1 | ln_1_land_144_lpi_1_dfm_1) & (~(ln_1_and_140_ssc_1
          | ln_1_land_146_lpi_1_dfm_1 | ln_1_land_147_lpi_1_dfm_1 | ln_1_land_148_lpi_1_dfm_1
          | ln_1_land_153_lpi_1_dfm_1 | ln_1_land_154_lpi_1_dfm_1 | ln_1_land_155_lpi_1_dfm_1
          | ln_1_land_156_lpi_1_dfm_1 | ln_1_land_161_lpi_1_dfm_1 | ln_1_land_162_lpi_1_dfm_1
          | ln_1_land_163_lpi_1_dfm_1 | ln_1_land_164_lpi_1_dfm_1 | ln_1_land_168_lpi_1_dfm_1
          | ln_1_land_169_lpi_1_dfm_1 | ln_1_land_170_lpi_1_dfm_1 | ln_1_land_171_lpi_1_dfm_1
          | ln_1_land_175_lpi_1_dfm_1 | ln_1_land_176_lpi_1_dfm_1 | ln_1_land_177_lpi_1_dfm_1
          | ln_1_land_181_lpi_1_dfm_1 | ln_1_land_182_lpi_1_dfm_1 | ln_1_land_183_lpi_1_dfm_1
          | ln_1_land_187_lpi_1_dfm_1 | ln_1_land_188_lpi_1_dfm_1 | ln_1_land_189_lpi_1_dfm_1
          | ln_1_land_193_lpi_1_dfm_1 | ln_1_land_194_lpi_1_dfm_1 | ln_1_land_198_lpi_1_dfm_1
          | ln_1_land_199_lpi_1_dfm_1 | ln_1_land_200_lpi_1_dfm_1 | ln_1_land_203_lpi_1_dfm_1
          | ln_1_land_204_lpi_1_dfm_1 | ln_1_land_208_lpi_1_dfm_1 | ln_1_land_209_lpi_1_dfm_1
          | ln_1_land_212_lpi_1_dfm_1 | ln_1_land_213_lpi_1_dfm_1 | ln_1_land_216_lpi_1_dfm_1
          | ln_1_land_217_lpi_1_dfm_1 | ln_1_land_220_lpi_1_dfm_1 | ln_1_land_221_lpi_1_dfm_1
          | ln_1_land_224_lpi_1_dfm_1 | ln_1_land_227_lpi_1_dfm_1 | ln_1_land_228_lpi_1_dfm_1
          | ln_1_land_230_lpi_1_dfm_1 | ln_1_land_231_lpi_1_dfm_1 | ln_1_land_233_lpi_1_dfm_1
          | ln_1_land_234_lpi_1_dfm_1 | ln_1_land_236_lpi_1_dfm_1 | ln_1_land_239_lpi_1_dfm_1
          | ln_1_land_241_lpi_1_dfm_1 | ln_1_land_243_lpi_1_dfm_1))) | ln_1_land_149_lpi_1_dfm_1
          | ln_1_land_150_lpi_1_dfm_1 | ln_1_land_151_lpi_1_dfm_1 | ln_1_land_152_lpi_1_dfm_1
          | ln_1_land_157_lpi_1_dfm_1 | ln_1_land_158_lpi_1_dfm_1 | ln_1_land_159_lpi_1_dfm_1
          | ln_1_land_160_lpi_1_dfm_1 | ln_1_land_165_lpi_1_dfm_1 | ln_1_land_166_lpi_1_dfm_1
          | ln_1_land_167_lpi_1_dfm_1 | ln_1_land_172_lpi_1_dfm_1 | ln_1_land_173_lpi_1_dfm_1
          | ln_1_land_174_lpi_1_dfm_1 | ln_1_land_178_lpi_1_dfm_1 | ln_1_land_179_lpi_1_dfm_1
          | ln_1_land_180_lpi_1_dfm_1 | ln_1_land_184_lpi_1_dfm_1 | ln_1_land_185_lpi_1_dfm_1
          | ln_1_land_186_lpi_1_dfm_1 | ln_1_land_190_lpi_1_dfm_1 | ln_1_land_191_lpi_1_dfm_1
          | ln_1_land_192_lpi_1_dfm_1 | ln_1_land_195_lpi_1_dfm_1 | ln_1_land_196_lpi_1_dfm_1
          | ln_1_land_197_lpi_1_dfm_1 | ln_1_land_201_lpi_1_dfm_1 | ln_1_land_202_lpi_1_dfm_1
          | ln_1_land_205_lpi_1_dfm_1 | ln_1_land_206_lpi_1_dfm_1 | ln_1_land_207_lpi_1_dfm_1
          | ln_1_land_210_lpi_1_dfm_1 | ln_1_land_211_lpi_1_dfm_1 | ln_1_land_214_lpi_1_dfm_1
          | ln_1_land_215_lpi_1_dfm_1 | ln_1_land_218_lpi_1_dfm_1 | ln_1_land_219_lpi_1_dfm_1
          | ln_1_land_222_lpi_1_dfm_1 | ln_1_land_223_lpi_1_dfm_1 | ln_1_land_225_lpi_1_dfm_1
          | ln_1_land_226_lpi_1_dfm_1 | ln_1_land_229_lpi_1_dfm_1 | ln_1_land_232_lpi_1_dfm_1
          | ln_1_land_235_lpi_1_dfm_1 | ln_1_land_237_lpi_1_dfm_1 | ln_1_land_238_lpi_1_dfm_1
          | ln_1_land_240_lpi_1_dfm_1 | ln_1_land_242_lpi_1_dfm_1 | ln_1_land_244_lpi_1_dfm_1;
      ln_1_ln_1_mux1h_118_psp_1_5 <= (((((~(((~(ln_1_ln_1_ln_1_nor_8_cse_1 | ln_1_land_6_lpi_1_dfm_1
          | ln_1_and_2_ssc_1)) & (~(ln_1_and_4_ssc_1 | ln_1_land_8_lpi_1_dfm_1 |
          ln_1_land_12_lpi_1_dfm_1 | ln_1_land_13_lpi_1_dfm_1 | ln_1_land_17_lpi_1_dfm_1
          | ln_1_land_18_lpi_1_dfm_1 | ln_1_land_21_lpi_1_dfm_1 | ln_1_land_22_lpi_1_dfm_1
          | ln_1_land_23_lpi_1_dfm_1 | ln_1_land_26_lpi_1_dfm_1 | ln_1_land_27_lpi_1_dfm_1
          | ln_1_land_30_lpi_1_dfm_1 | ln_1_land_31_lpi_1_dfm_1 | ln_1_land_35_lpi_1_dfm_1
          | ln_1_land_36_lpi_1_dfm_1 | ln_1_land_39_lpi_1_dfm_1 | ln_1_land_40_lpi_1_dfm_1
          | ln_1_land_43_lpi_1_dfm_1 | ln_1_land_44_lpi_1_dfm_1 | ln_1_land_47_lpi_1_dfm_1
          | ln_1_land_48_lpi_1_dfm_1))) | ln_1_land_9_lpi_1_dfm_1 | ln_1_land_10_lpi_1_dfm_1
          | ln_1_land_11_lpi_1_dfm_1 | ln_1_land_14_lpi_1_dfm_1 | ln_1_land_15_lpi_1_dfm_1
          | ln_1_land_16_lpi_1_dfm_1 | ln_1_land_19_lpi_1_dfm_1 | ln_1_land_20_lpi_1_dfm_1
          | ln_1_land_24_lpi_1_dfm_1 | ln_1_land_25_lpi_1_dfm_1 | ln_1_land_28_lpi_1_dfm_1
          | ln_1_land_29_lpi_1_dfm_1 | ln_1_land_32_lpi_1_dfm_1 | ln_1_land_33_lpi_1_dfm_1
          | ln_1_land_34_lpi_1_dfm_1 | ln_1_land_37_lpi_1_dfm_1 | ln_1_land_38_lpi_1_dfm_1
          | ln_1_land_41_lpi_1_dfm_1 | ln_1_land_42_lpi_1_dfm_1 | ln_1_land_45_lpi_1_dfm_1
          | ln_1_land_46_lpi_1_dfm_1 | ln_1_land_49_lpi_1_dfm_1 | ln_1_if_50_ln_1_if_50_and_seb_1
          | ln_1_land_52_lpi_1_dfm_1)) | ln_1_land_51_lpi_1_dfm_1) & (~(ln_1_and_48_ssc_1
          | ln_1_land_56_lpi_1_dfm_1 | ln_1_land_57_lpi_1_dfm_1 | ln_1_land_60_lpi_1_dfm_1
          | ln_1_land_63_lpi_1_dfm_1 | ln_1_land_64_lpi_1_dfm_1 | ln_1_land_66_lpi_1_dfm_1
          | ln_1_land_67_lpi_1_dfm_1 | ln_1_land_69_lpi_1_dfm_1 | ln_1_land_70_lpi_1_dfm_1
          | ln_1_land_73_lpi_1_dfm_1 | ln_1_land_76_lpi_1_dfm_1 | ln_1_land_79_lpi_1_dfm_1
          | ln_1_land_81_lpi_1_dfm_1 | ln_1_land_82_lpi_1_dfm_1 | ln_1_land_84_lpi_1_dfm_1
          | ln_1_land_87_lpi_1_dfm_1 | ln_1_land_89_lpi_1_dfm_1 | ln_1_land_90_lpi_1_dfm_1
          | ln_1_land_92_lpi_1_dfm_1 | ln_1_land_94_lpi_1_dfm_1 | ln_1_land_97_lpi_1_dfm_1
          | ln_1_land_99_lpi_1_dfm_1 | ln_1_land_101_lpi_1_dfm_1 | ln_1_land_103_lpi_1_dfm_1
          | ln_1_land_105_lpi_1_dfm_1 | ln_1_land_107_lpi_1_dfm_1 | ln_1_land_109_lpi_1_dfm_1
          | ln_1_land_111_lpi_1_dfm_1 | ln_1_land_113_lpi_1_dfm_1 | ln_1_land_115_lpi_1_dfm_1
          | ln_1_land_116_lpi_1_dfm_1 | ln_1_land_118_lpi_1_dfm_1 | ln_1_land_120_lpi_1_dfm_1
          | ln_1_land_121_lpi_1_dfm_1 | ln_1_land_125_lpi_1_dfm_1 | ln_1_land_126_lpi_1_dfm_1
          | ln_1_land_130_lpi_1_dfm_1 | ln_1_land_131_lpi_1_dfm_1 | ln_1_land_134_lpi_1_dfm_1
          | ln_1_land_135_lpi_1_dfm_1 | ln_1_land_136_lpi_1_dfm_1 | ln_1_land_139_lpi_1_dfm_1
          | ln_1_land_140_lpi_1_dfm_1))) | ln_1_land_54_lpi_1_dfm_1 | ln_1_land_55_lpi_1_dfm_1
          | ln_1_land_58_lpi_1_dfm_1 | ln_1_land_59_lpi_1_dfm_1 | ln_1_land_61_lpi_1_dfm_1
          | ln_1_land_62_lpi_1_dfm_1 | ln_1_land_65_lpi_1_dfm_1 | ln_1_land_68_lpi_1_dfm_1
          | ln_1_land_71_lpi_1_dfm_1 | ln_1_land_72_lpi_1_dfm_1 | ln_1_land_74_lpi_1_dfm_1
          | ln_1_land_75_lpi_1_dfm_1 | ln_1_land_77_lpi_1_dfm_1 | ln_1_land_78_lpi_1_dfm_1
          | ln_1_land_80_lpi_1_dfm_1 | ln_1_land_83_lpi_1_dfm_1 | ln_1_land_85_lpi_1_dfm_1
          | ln_1_land_86_lpi_1_dfm_1 | ln_1_land_88_lpi_1_dfm_1 | ln_1_land_91_lpi_1_dfm_1
          | ln_1_land_93_lpi_1_dfm_1 | ln_1_land_95_lpi_1_dfm_1 | ln_1_land_96_lpi_1_dfm_1
          | ln_1_land_98_lpi_1_dfm_1 | ln_1_land_100_lpi_1_dfm_1 | ln_1_land_102_lpi_1_dfm_1
          | ln_1_land_104_lpi_1_dfm_1 | ln_1_land_106_lpi_1_dfm_1 | ln_1_land_108_lpi_1_dfm_1
          | ln_1_land_110_lpi_1_dfm_1 | ln_1_land_112_lpi_1_dfm_1 | ln_1_land_114_lpi_1_dfm_1
          | ln_1_land_117_lpi_1_dfm_1 | ln_1_land_119_lpi_1_dfm_1 | ln_1_land_122_lpi_1_dfm_1
          | ln_1_land_123_lpi_1_dfm_1 | ln_1_land_124_lpi_1_dfm_1 | ln_1_land_127_lpi_1_dfm_1
          | ln_1_land_128_lpi_1_dfm_1 | ln_1_land_129_lpi_1_dfm_1 | ln_1_land_132_lpi_1_dfm_1
          | ln_1_land_133_lpi_1_dfm_1 | ln_1_land_137_lpi_1_dfm_1 | ln_1_land_138_lpi_1_dfm_1
          | ln_1_land_141_lpi_1_dfm_1 | ln_1_land_142_lpi_1_dfm_1) & ln_1_nor_3_cse_1
          & (~(ln_1_land_147_lpi_1_dfm_1 | ln_1_land_148_lpi_1_dfm_1 | ln_1_land_151_lpi_1_dfm_1
          | ln_1_land_152_lpi_1_dfm_1 | ln_1_land_155_lpi_1_dfm_1 | ln_1_land_156_lpi_1_dfm_1
          | ln_1_land_159_lpi_1_dfm_1 | ln_1_land_160_lpi_1_dfm_1 | ln_1_land_163_lpi_1_dfm_1
          | ln_1_land_164_lpi_1_dfm_1 | ln_1_land_166_lpi_1_dfm_1 | ln_1_land_167_lpi_1_dfm_1
          | ln_1_land_170_lpi_1_dfm_1 | ln_1_land_171_lpi_1_dfm_1 | ln_1_land_173_lpi_1_dfm_1
          | ln_1_land_174_lpi_1_dfm_1 | ln_1_land_177_lpi_1_dfm_1 | ln_1_land_180_lpi_1_dfm_1
          | ln_1_land_183_lpi_1_dfm_1 | ln_1_land_186_lpi_1_dfm_1 | ln_1_land_189_lpi_1_dfm_1
          | ln_1_land_191_lpi_1_dfm_1 | ln_1_land_192_lpi_1_dfm_1 | ln_1_land_194_lpi_1_dfm_1
          | ln_1_land_197_lpi_1_dfm_1 | ln_1_land_199_lpi_1_dfm_1 | ln_1_land_200_lpi_1_dfm_1
          | ln_1_land_202_lpi_1_dfm_1 | ln_1_land_204_lpi_1_dfm_1 | ln_1_land_206_lpi_1_dfm_1
          | ln_1_land_207_lpi_1_dfm_1 | ln_1_land_209_lpi_1_dfm_1 | ln_1_land_211_lpi_1_dfm_1
          | ln_1_land_213_lpi_1_dfm_1 | ln_1_land_215_lpi_1_dfm_1 | ln_1_land_217_lpi_1_dfm_1
          | ln_1_land_219_lpi_1_dfm_1 | ln_1_land_221_lpi_1_dfm_1 | ln_1_land_223_lpi_1_dfm_1
          | ln_1_land_224_lpi_1_dfm_1 | ln_1_land_226_lpi_1_dfm_1 | ln_1_land_228_lpi_1_dfm_1
          | ln_1_land_229_lpi_1_dfm_1 | ln_1_land_231_lpi_1_dfm_1 | ln_1_land_232_lpi_1_dfm_1
          | ln_1_land_234_lpi_1_dfm_1 | ln_1_land_235_lpi_1_dfm_1 | ln_1_land_238_lpi_1_dfm_1
          | ln_1_land_239_lpi_1_dfm_1 | ln_1_land_240_lpi_1_dfm_1))) | ln_1_and_140_ssc_1
          | ln_1_land_146_lpi_1_dfm_1 | ln_1_land_149_lpi_1_dfm_1 | ln_1_land_150_lpi_1_dfm_1
          | ln_1_land_153_lpi_1_dfm_1 | ln_1_land_154_lpi_1_dfm_1 | ln_1_land_157_lpi_1_dfm_1
          | ln_1_land_158_lpi_1_dfm_1 | ln_1_land_161_lpi_1_dfm_1 | ln_1_land_162_lpi_1_dfm_1
          | ln_1_land_165_lpi_1_dfm_1 | ln_1_land_168_lpi_1_dfm_1 | ln_1_land_169_lpi_1_dfm_1
          | ln_1_land_172_lpi_1_dfm_1 | ln_1_land_175_lpi_1_dfm_1 | ln_1_land_176_lpi_1_dfm_1
          | ln_1_land_178_lpi_1_dfm_1 | ln_1_land_179_lpi_1_dfm_1 | ln_1_land_181_lpi_1_dfm_1
          | ln_1_land_182_lpi_1_dfm_1 | ln_1_land_184_lpi_1_dfm_1 | ln_1_land_185_lpi_1_dfm_1
          | ln_1_land_187_lpi_1_dfm_1 | ln_1_land_188_lpi_1_dfm_1 | ln_1_land_190_lpi_1_dfm_1
          | ln_1_land_193_lpi_1_dfm_1 | ln_1_land_195_lpi_1_dfm_1 | ln_1_land_196_lpi_1_dfm_1
          | ln_1_land_198_lpi_1_dfm_1 | ln_1_land_201_lpi_1_dfm_1 | ln_1_land_203_lpi_1_dfm_1
          | ln_1_land_205_lpi_1_dfm_1 | ln_1_land_208_lpi_1_dfm_1 | ln_1_land_210_lpi_1_dfm_1
          | ln_1_land_212_lpi_1_dfm_1 | ln_1_land_214_lpi_1_dfm_1 | ln_1_land_216_lpi_1_dfm_1
          | ln_1_land_218_lpi_1_dfm_1 | ln_1_land_220_lpi_1_dfm_1 | ln_1_land_222_lpi_1_dfm_1
          | ln_1_land_225_lpi_1_dfm_1 | ln_1_land_227_lpi_1_dfm_1 | ln_1_land_230_lpi_1_dfm_1
          | ln_1_land_233_lpi_1_dfm_1 | ln_1_land_236_lpi_1_dfm_1 | ln_1_land_237_lpi_1_dfm_1
          | ln_1_land_241_lpi_1_dfm_1 | ln_1_land_242_lpi_1_dfm_1 | ln_1_land_243_lpi_1_dfm_1
          | ln_1_land_244_lpi_1_dfm_1;
      ln_1_ln_1_mux1h_118_psp_1_4 <= (((~((~((~((~((((~(((~((~((~(ln_1_ret_13_0_lpi_1_dfm_257
          | ln_1_land_3_lpi_1_dfm_1)) | ln_1_land_4_lpi_1_dfm_1 | ln_1_land_6_lpi_1_dfm_1))
          | ln_1_and_2_ssc_1)) & (~(ln_1_and_4_ssc_1 | ln_1_land_9_lpi_1_dfm_1 |
          ln_1_land_12_lpi_1_dfm_1 | ln_1_land_14_lpi_1_dfm_1 | ln_1_land_17_lpi_1_dfm_1
          | ln_1_land_19_lpi_1_dfm_1 | ln_1_land_21_lpi_1_dfm_1 | ln_1_land_24_lpi_1_dfm_1
          | ln_1_land_26_lpi_1_dfm_1 | ln_1_land_28_lpi_1_dfm_1 | ln_1_land_30_lpi_1_dfm_1
          | ln_1_land_32_lpi_1_dfm_1 | ln_1_land_33_lpi_1_dfm_1 | ln_1_land_35_lpi_1_dfm_1
          | ln_1_land_37_lpi_1_dfm_1 | ln_1_land_39_lpi_1_dfm_1 | ln_1_land_41_lpi_1_dfm_1
          | ln_1_land_43_lpi_1_dfm_1 | ln_1_land_45_lpi_1_dfm_1 | ln_1_land_47_lpi_1_dfm_1
          | ln_1_land_49_lpi_1_dfm_1))) | ln_1_land_8_lpi_1_dfm_1 | ln_1_land_10_lpi_1_dfm_1
          | ln_1_land_11_lpi_1_dfm_1 | ln_1_land_13_lpi_1_dfm_1 | ln_1_land_15_lpi_1_dfm_1
          | ln_1_land_16_lpi_1_dfm_1 | ln_1_land_18_lpi_1_dfm_1 | ln_1_land_20_lpi_1_dfm_1
          | ln_1_land_22_lpi_1_dfm_1 | ln_1_land_23_lpi_1_dfm_1 | ln_1_land_25_lpi_1_dfm_1
          | ln_1_land_27_lpi_1_dfm_1 | ln_1_land_29_lpi_1_dfm_1 | ln_1_land_31_lpi_1_dfm_1
          | ln_1_land_34_lpi_1_dfm_1 | ln_1_land_36_lpi_1_dfm_1 | ln_1_land_38_lpi_1_dfm_1
          | ln_1_land_40_lpi_1_dfm_1 | ln_1_land_42_lpi_1_dfm_1 | ln_1_land_44_lpi_1_dfm_1
          | ln_1_land_46_lpi_1_dfm_1 | ln_1_land_48_lpi_1_dfm_1 | ln_1_if_50_ln_1_if_50_and_seb_1
          | ln_1_land_51_lpi_1_dfm_1)) | ln_1_land_52_lpi_1_dfm_1) & (~(ln_1_and_48_ssc_1
          | ln_1_land_55_lpi_1_dfm_1 | ln_1_land_57_lpi_1_dfm_1 | ln_1_land_59_lpi_1_dfm_1
          | ln_1_land_60_lpi_1_dfm_1 | ln_1_land_62_lpi_1_dfm_1 | ln_1_land_64_lpi_1_dfm_1
          | ln_1_land_65_lpi_1_dfm_1 | ln_1_land_67_lpi_1_dfm_1 | ln_1_land_70_lpi_1_dfm_1
          | ln_1_land_72_lpi_1_dfm_1 | ln_1_land_73_lpi_1_dfm_1 | ln_1_land_75_lpi_1_dfm_1
          | ln_1_land_76_lpi_1_dfm_1 | ln_1_land_78_lpi_1_dfm_1 | ln_1_land_79_lpi_1_dfm_1
          | ln_1_land_82_lpi_1_dfm_1 | ln_1_land_83_lpi_1_dfm_1 | ln_1_land_86_lpi_1_dfm_1
          | ln_1_land_87_lpi_1_dfm_1 | ln_1_land_90_lpi_1_dfm_1 | ln_1_land_91_lpi_1_dfm_1
          | ln_1_land_92_lpi_1_dfm_1 | ln_1_land_96_lpi_1_dfm_1 | ln_1_land_97_lpi_1_dfm_1
          | ln_1_land_98_lpi_1_dfm_1 | ln_1_land_99_lpi_1_dfm_1 | ln_1_land_100_lpi_1_dfm_1
          | ln_1_land_112_lpi_1_dfm_1 | ln_1_land_113_lpi_1_dfm_1 | ln_1_land_114_lpi_1_dfm_1
          | ln_1_land_115_lpi_1_dfm_1 | ln_1_land_118_lpi_1_dfm_1 | ln_1_land_119_lpi_1_dfm_1
          | ln_1_land_121_lpi_1_dfm_1 | ln_1_land_124_lpi_1_dfm_1 | ln_1_land_126_lpi_1_dfm_1
          | ln_1_land_128_lpi_1_dfm_1 | ln_1_land_129_lpi_1_dfm_1 | ln_1_land_131_lpi_1_dfm_1
          | ln_1_land_133_lpi_1_dfm_1 | ln_1_land_135_lpi_1_dfm_1 | ln_1_land_136_lpi_1_dfm_1
          | ln_1_land_138_lpi_1_dfm_1 | ln_1_land_140_lpi_1_dfm_1))) | ln_1_land_54_lpi_1_dfm_1
          | ln_1_land_56_lpi_1_dfm_1 | ln_1_land_58_lpi_1_dfm_1 | ln_1_land_61_lpi_1_dfm_1
          | ln_1_land_63_lpi_1_dfm_1 | ln_1_land_66_lpi_1_dfm_1 | ln_1_land_68_lpi_1_dfm_1
          | ln_1_land_69_lpi_1_dfm_1 | ln_1_land_71_lpi_1_dfm_1 | ln_1_land_74_lpi_1_dfm_1
          | ln_1_land_77_lpi_1_dfm_1 | ln_1_land_80_lpi_1_dfm_1 | ln_1_land_81_lpi_1_dfm_1
          | ln_1_land_84_lpi_1_dfm_1 | ln_1_land_85_lpi_1_dfm_1 | ln_1_land_88_lpi_1_dfm_1
          | ln_1_land_89_lpi_1_dfm_1 | ln_1_land_93_lpi_1_dfm_1 | ln_1_land_94_lpi_1_dfm_1
          | ln_1_land_95_lpi_1_dfm_1 | ln_1_land_101_lpi_1_dfm_1 | ln_1_land_102_lpi_1_dfm_1
          | ln_1_land_103_lpi_1_dfm_1 | ln_1_land_104_lpi_1_dfm_1 | ln_1_land_105_lpi_1_dfm_1
          | ln_1_land_106_lpi_1_dfm_1 | ln_1_land_107_lpi_1_dfm_1 | ln_1_land_108_lpi_1_dfm_1
          | ln_1_land_109_lpi_1_dfm_1 | ln_1_land_110_lpi_1_dfm_1 | ln_1_land_111_lpi_1_dfm_1
          | ln_1_land_116_lpi_1_dfm_1 | ln_1_land_117_lpi_1_dfm_1 | ln_1_land_120_lpi_1_dfm_1
          | ln_1_land_122_lpi_1_dfm_1 | ln_1_land_123_lpi_1_dfm_1 | ln_1_land_125_lpi_1_dfm_1
          | ln_1_land_127_lpi_1_dfm_1 | ln_1_land_130_lpi_1_dfm_1 | ln_1_land_132_lpi_1_dfm_1
          | ln_1_land_134_lpi_1_dfm_1 | ln_1_land_137_lpi_1_dfm_1 | ln_1_land_139_lpi_1_dfm_1))
          | ln_1_land_142_lpi_1_dfm_1)) | ln_1_land_141_lpi_1_dfm_1)) | ln_1_land_144_lpi_1_dfm_1))
          | ln_1_and_138_ssc_1) & (~(ln_1_land_146_lpi_1_dfm_1 | ln_1_land_148_lpi_1_dfm_1
          | ln_1_land_150_lpi_1_dfm_1 | ln_1_land_152_lpi_1_dfm_1 | ln_1_land_154_lpi_1_dfm_1
          | ln_1_land_156_lpi_1_dfm_1 | ln_1_land_158_lpi_1_dfm_1 | ln_1_land_160_lpi_1_dfm_1
          | ln_1_land_162_lpi_1_dfm_1 | ln_1_land_164_lpi_1_dfm_1 | ln_1_land_167_lpi_1_dfm_1
          | ln_1_land_169_lpi_1_dfm_1 | ln_1_land_171_lpi_1_dfm_1 | ln_1_land_172_lpi_1_dfm_1
          | ln_1_land_174_lpi_1_dfm_1 | ln_1_land_176_lpi_1_dfm_1 | ln_1_land_177_lpi_1_dfm_1
          | ln_1_land_179_lpi_1_dfm_1 | ln_1_land_180_lpi_1_dfm_1 | ln_1_land_182_lpi_1_dfm_1
          | ln_1_land_185_lpi_1_dfm_1 | ln_1_land_186_lpi_1_dfm_1 | ln_1_land_188_lpi_1_dfm_1
          | ln_1_land_189_lpi_1_dfm_1 | ln_1_land_192_lpi_1_dfm_1 | ln_1_land_193_lpi_1_dfm_1
          | ln_1_land_196_lpi_1_dfm_1 | ln_1_land_197_lpi_1_dfm_1 | ln_1_land_200_lpi_1_dfm_1
          | ln_1_land_201_lpi_1_dfm_1 | ln_1_land_202_lpi_1_dfm_1 | ln_1_land_207_lpi_1_dfm_1
          | ln_1_land_208_lpi_1_dfm_1 | ln_1_land_209_lpi_1_dfm_1 | ln_1_land_210_lpi_1_dfm_1
          | ln_1_land_211_lpi_1_dfm_1 | ln_1_land_212_lpi_1_dfm_1 | ln_1_land_218_lpi_1_dfm_1
          | ln_1_land_219_lpi_1_dfm_1 | ln_1_land_220_lpi_1_dfm_1 | ln_1_land_221_lpi_1_dfm_1
          | ln_1_land_222_lpi_1_dfm_1 | ln_1_land_223_lpi_1_dfm_1 | ln_1_land_226_lpi_1_dfm_1
          | ln_1_land_227_lpi_1_dfm_1 | ln_1_land_228_lpi_1_dfm_1 | ln_1_land_230_lpi_1_dfm_1
          | ln_1_land_231_lpi_1_dfm_1 | ln_1_land_233_lpi_1_dfm_1 | ln_1_land_234_lpi_1_dfm_1
          | ln_1_land_236_lpi_1_dfm_1 | ln_1_land_238_lpi_1_dfm_1 | ln_1_land_239_lpi_1_dfm_1
          | ln_1_land_241_lpi_1_dfm_1 | ln_1_land_242_lpi_1_dfm_1))) | ln_1_and_140_ssc_1
          | ln_1_land_147_lpi_1_dfm_1 | ln_1_land_149_lpi_1_dfm_1 | ln_1_land_151_lpi_1_dfm_1
          | ln_1_land_153_lpi_1_dfm_1 | ln_1_land_155_lpi_1_dfm_1 | ln_1_land_157_lpi_1_dfm_1
          | ln_1_land_159_lpi_1_dfm_1 | ln_1_land_161_lpi_1_dfm_1 | ln_1_land_163_lpi_1_dfm_1
          | ln_1_land_165_lpi_1_dfm_1 | ln_1_land_166_lpi_1_dfm_1 | ln_1_land_168_lpi_1_dfm_1
          | ln_1_land_170_lpi_1_dfm_1 | ln_1_land_173_lpi_1_dfm_1 | ln_1_land_175_lpi_1_dfm_1
          | ln_1_land_178_lpi_1_dfm_1 | ln_1_land_181_lpi_1_dfm_1 | ln_1_land_183_lpi_1_dfm_1
          | ln_1_land_184_lpi_1_dfm_1 | ln_1_land_187_lpi_1_dfm_1 | ln_1_land_190_lpi_1_dfm_1
          | ln_1_land_191_lpi_1_dfm_1 | ln_1_land_194_lpi_1_dfm_1 | ln_1_land_195_lpi_1_dfm_1
          | ln_1_land_198_lpi_1_dfm_1 | ln_1_land_199_lpi_1_dfm_1 | ln_1_land_203_lpi_1_dfm_1
          | ln_1_land_204_lpi_1_dfm_1 | ln_1_land_205_lpi_1_dfm_1 | ln_1_land_206_lpi_1_dfm_1
          | ln_1_land_213_lpi_1_dfm_1 | ln_1_land_214_lpi_1_dfm_1 | ln_1_land_215_lpi_1_dfm_1
          | ln_1_land_216_lpi_1_dfm_1 | ln_1_land_217_lpi_1_dfm_1 | ln_1_land_224_lpi_1_dfm_1
          | ln_1_land_225_lpi_1_dfm_1 | ln_1_land_229_lpi_1_dfm_1 | ln_1_land_232_lpi_1_dfm_1
          | ln_1_land_235_lpi_1_dfm_1 | ln_1_land_237_lpi_1_dfm_1 | ln_1_land_240_lpi_1_dfm_1
          | ln_1_land_243_lpi_1_dfm_1 | ln_1_land_244_lpi_1_dfm_1;
      ln_1_ln_1_mux1h_118_psp_1_3 <= (((~((~((((~(((~((~(ln_1_ret_13_0_lpi_1_dfm_257
          | ln_1_land_3_lpi_1_dfm_1 | ln_1_land_4_lpi_1_dfm_1 | ln_1_land_6_lpi_1_dfm_1))
          | ln_1_and_2_ssc_1)) & (~(ln_1_land_9_lpi_1_dfm_1 | ln_1_land_10_lpi_1_dfm_1
          | ln_1_land_14_lpi_1_dfm_1 | ln_1_land_15_lpi_1_dfm_1 | ln_1_land_20_lpi_1_dfm_1
          | ln_1_land_21_lpi_1_dfm_1 | ln_1_land_22_lpi_1_dfm_1 | ln_1_land_27_lpi_1_dfm_1
          | ln_1_land_28_lpi_1_dfm_1 | ln_1_land_29_lpi_1_dfm_1 | ln_1_land_30_lpi_1_dfm_1
          | ln_1_land_31_lpi_1_dfm_1 | ln_1_land_32_lpi_1_dfm_1))) | ln_1_and_4_ssc_1
          | ln_1_land_8_lpi_1_dfm_1 | ln_1_land_11_lpi_1_dfm_1 | ln_1_land_12_lpi_1_dfm_1
          | ln_1_land_13_lpi_1_dfm_1 | ln_1_land_16_lpi_1_dfm_1 | ln_1_land_17_lpi_1_dfm_1
          | ln_1_land_18_lpi_1_dfm_1 | ln_1_land_19_lpi_1_dfm_1 | ln_1_land_23_lpi_1_dfm_1
          | ln_1_land_24_lpi_1_dfm_1 | ln_1_land_25_lpi_1_dfm_1 | ln_1_land_26_lpi_1_dfm_1
          | ln_1_land_33_lpi_1_dfm_1 | ln_1_land_34_lpi_1_dfm_1 | ln_1_land_35_lpi_1_dfm_1
          | ln_1_land_36_lpi_1_dfm_1 | ln_1_land_37_lpi_1_dfm_1 | ln_1_land_38_lpi_1_dfm_1
          | ln_1_land_39_lpi_1_dfm_1 | ln_1_land_40_lpi_1_dfm_1 | ln_1_land_41_lpi_1_dfm_1
          | ln_1_land_42_lpi_1_dfm_1 | ln_1_land_43_lpi_1_dfm_1 | ln_1_land_44_lpi_1_dfm_1
          | ln_1_land_45_lpi_1_dfm_1 | ln_1_land_46_lpi_1_dfm_1 | ln_1_land_47_lpi_1_dfm_1
          | ln_1_land_48_lpi_1_dfm_1 | ln_1_land_49_lpi_1_dfm_1 | ln_1_if_50_ln_1_if_50_and_seb_1))
          | ln_1_land_51_lpi_1_dfm_1 | ln_1_land_52_lpi_1_dfm_1) & (~(ln_1_land_56_lpi_1_dfm_1
          | ln_1_land_57_lpi_1_dfm_1 | ln_1_land_58_lpi_1_dfm_1 | ln_1_land_59_lpi_1_dfm_1
          | ln_1_land_63_lpi_1_dfm_1 | ln_1_land_64_lpi_1_dfm_1 | ln_1_land_67_lpi_1_dfm_1
          | ln_1_land_68_lpi_1_dfm_1 | ln_1_land_71_lpi_1_dfm_1 | ln_1_land_72_lpi_1_dfm_1
          | ln_1_land_74_lpi_1_dfm_1 | ln_1_land_75_lpi_1_dfm_1 | ln_1_land_77_lpi_1_dfm_1
          | ln_1_land_78_lpi_1_dfm_1 | ln_1_land_80_lpi_1_dfm_1 | ln_1_land_82_lpi_1_dfm_1
          | ln_1_land_84_lpi_1_dfm_1 | ln_1_land_86_lpi_1_dfm_1 | ln_1_land_88_lpi_1_dfm_1
          | ln_1_land_90_lpi_1_dfm_1 | ln_1_land_91_lpi_1_dfm_1 | ln_1_land_93_lpi_1_dfm_1
          | ln_1_land_96_lpi_1_dfm_1 | ln_1_land_97_lpi_1_dfm_1 | ln_1_land_101_lpi_1_dfm_1
          | ln_1_land_102_lpi_1_dfm_1 | ln_1_land_103_lpi_1_dfm_1 | ln_1_land_104_lpi_1_dfm_1
          | ln_1_land_105_lpi_1_dfm_1 | ln_1_land_107_lpi_1_dfm_1 | ln_1_land_108_lpi_1_dfm_1
          | ln_1_land_109_lpi_1_dfm_1 | ln_1_land_110_lpi_1_dfm_1 | ln_1_land_111_lpi_1_dfm_1
          | ln_1_land_114_lpi_1_dfm_1 | ln_1_land_115_lpi_1_dfm_1 | ln_1_land_117_lpi_1_dfm_1
          | ln_1_land_119_lpi_1_dfm_1 | ln_1_land_123_lpi_1_dfm_1 | ln_1_land_124_lpi_1_dfm_1
          | ln_1_land_129_lpi_1_dfm_1 | ln_1_land_130_lpi_1_dfm_1 | ln_1_land_131_lpi_1_dfm_1
          | ln_1_land_136_lpi_1_dfm_1 | ln_1_land_137_lpi_1_dfm_1 | ln_1_land_138_lpi_1_dfm_1
          | ln_1_land_139_lpi_1_dfm_1 | ln_1_land_140_lpi_1_dfm_1))) | ln_1_and_48_ssc_1
          | ln_1_land_54_lpi_1_dfm_1 | ln_1_land_55_lpi_1_dfm_1 | ln_1_land_60_lpi_1_dfm_1
          | ln_1_land_61_lpi_1_dfm_1 | ln_1_land_62_lpi_1_dfm_1 | ln_1_land_65_lpi_1_dfm_1
          | ln_1_land_66_lpi_1_dfm_1 | ln_1_land_69_lpi_1_dfm_1 | ln_1_land_70_lpi_1_dfm_1
          | ln_1_land_73_lpi_1_dfm_1 | ln_1_land_76_lpi_1_dfm_1 | ln_1_land_79_lpi_1_dfm_1
          | ln_1_land_81_lpi_1_dfm_1 | ln_1_land_83_lpi_1_dfm_1 | ln_1_land_85_lpi_1_dfm_1
          | ln_1_land_87_lpi_1_dfm_1 | ln_1_land_89_lpi_1_dfm_1 | ln_1_land_92_lpi_1_dfm_1
          | ln_1_land_94_lpi_1_dfm_1 | ln_1_land_95_lpi_1_dfm_1 | ln_1_land_98_lpi_1_dfm_1
          | ln_1_land_99_lpi_1_dfm_1 | ln_1_land_100_lpi_1_dfm_1 | ln_1_land_106_lpi_1_dfm_1
          | ln_1_land_112_lpi_1_dfm_1 | ln_1_land_113_lpi_1_dfm_1 | ln_1_land_116_lpi_1_dfm_1
          | ln_1_land_118_lpi_1_dfm_1 | ln_1_land_120_lpi_1_dfm_1 | ln_1_land_121_lpi_1_dfm_1
          | ln_1_land_122_lpi_1_dfm_1 | ln_1_land_125_lpi_1_dfm_1 | ln_1_land_126_lpi_1_dfm_1
          | ln_1_land_127_lpi_1_dfm_1 | ln_1_land_128_lpi_1_dfm_1 | ln_1_land_132_lpi_1_dfm_1
          | ln_1_land_133_lpi_1_dfm_1 | ln_1_land_134_lpi_1_dfm_1 | ln_1_land_135_lpi_1_dfm_1))
          | ln_1_land_141_lpi_1_dfm_1)) | ln_1_land_142_lpi_1_dfm_1 | ln_1_and_138_ssc_1
          | ln_1_land_144_lpi_1_dfm_1) & (~(ln_1_land_160_lpi_1_dfm_1 | ln_1_land_161_lpi_1_dfm_1
          | ln_1_land_162_lpi_1_dfm_1 | ln_1_land_163_lpi_1_dfm_1 | ln_1_land_164_lpi_1_dfm_1
          | ln_1_land_165_lpi_1_dfm_1 | ln_1_land_169_lpi_1_dfm_1 | ln_1_land_170_lpi_1_dfm_1
          | ln_1_land_171_lpi_1_dfm_1 | ln_1_land_174_lpi_1_dfm_1 | ln_1_land_175_lpi_1_dfm_1
          | ln_1_land_176_lpi_1_dfm_1 | ln_1_land_179_lpi_1_dfm_1 | ln_1_land_182_lpi_1_dfm_1
          | ln_1_land_183_lpi_1_dfm_1 | ln_1_land_185_lpi_1_dfm_1 | ln_1_land_188_lpi_1_dfm_1
          | ln_1_land_190_lpi_1_dfm_1 | ln_1_land_192_lpi_1_dfm_1 | ln_1_land_194_lpi_1_dfm_1
          | ln_1_land_196_lpi_1_dfm_1 | ln_1_land_198_lpi_1_dfm_1 | ln_1_land_200_lpi_1_dfm_1
          | ln_1_land_201_lpi_1_dfm_1 | ln_1_land_203_lpi_1_dfm_1 | ln_1_land_204_lpi_1_dfm_1
          | ln_1_land_207_lpi_1_dfm_1 | ln_1_land_208_lpi_1_dfm_1 | ln_1_land_213_lpi_1_dfm_1
          | ln_1_land_214_lpi_1_dfm_1 | ln_1_land_215_lpi_1_dfm_1 | ln_1_land_216_lpi_1_dfm_1
          | ln_1_land_217_lpi_1_dfm_1 | ln_1_land_222_lpi_1_dfm_1 | ln_1_land_223_lpi_1_dfm_1
          | ln_1_land_225_lpi_1_dfm_1 | ln_1_land_228_lpi_1_dfm_1 | ln_1_land_231_lpi_1_dfm_1
          | ln_1_land_234_lpi_1_dfm_1 | ln_1_land_235_lpi_1_dfm_1 | ln_1_land_236_lpi_1_dfm_1
          | ln_1_land_237_lpi_1_dfm_1 | ln_1_land_238_lpi_1_dfm_1 | ln_1_land_241_lpi_1_dfm_1
          | ln_1_land_243_lpi_1_dfm_1))) | ln_1_and_140_ssc_1 | ln_1_land_146_lpi_1_dfm_1
          | ln_1_land_147_lpi_1_dfm_1 | ln_1_land_148_lpi_1_dfm_1 | ln_1_land_149_lpi_1_dfm_1
          | ln_1_land_150_lpi_1_dfm_1 | ln_1_land_151_lpi_1_dfm_1 | ln_1_land_152_lpi_1_dfm_1
          | ln_1_land_153_lpi_1_dfm_1 | ln_1_land_154_lpi_1_dfm_1 | ln_1_land_155_lpi_1_dfm_1
          | ln_1_land_156_lpi_1_dfm_1 | ln_1_land_157_lpi_1_dfm_1 | ln_1_land_158_lpi_1_dfm_1
          | ln_1_land_159_lpi_1_dfm_1 | ln_1_land_166_lpi_1_dfm_1 | ln_1_land_167_lpi_1_dfm_1
          | ln_1_land_168_lpi_1_dfm_1 | ln_1_land_172_lpi_1_dfm_1 | ln_1_land_173_lpi_1_dfm_1
          | ln_1_land_177_lpi_1_dfm_1 | ln_1_land_178_lpi_1_dfm_1 | ln_1_land_180_lpi_1_dfm_1
          | ln_1_land_181_lpi_1_dfm_1 | ln_1_land_184_lpi_1_dfm_1 | ln_1_land_186_lpi_1_dfm_1
          | ln_1_land_187_lpi_1_dfm_1 | ln_1_land_189_lpi_1_dfm_1 | ln_1_land_191_lpi_1_dfm_1
          | ln_1_land_193_lpi_1_dfm_1 | ln_1_land_195_lpi_1_dfm_1 | ln_1_land_197_lpi_1_dfm_1
          | ln_1_land_199_lpi_1_dfm_1 | ln_1_land_202_lpi_1_dfm_1 | ln_1_land_205_lpi_1_dfm_1
          | ln_1_land_206_lpi_1_dfm_1 | ln_1_land_209_lpi_1_dfm_1 | ln_1_land_210_lpi_1_dfm_1
          | ln_1_land_211_lpi_1_dfm_1 | ln_1_land_212_lpi_1_dfm_1 | ln_1_land_218_lpi_1_dfm_1
          | ln_1_land_219_lpi_1_dfm_1 | ln_1_land_220_lpi_1_dfm_1 | ln_1_land_221_lpi_1_dfm_1
          | ln_1_land_224_lpi_1_dfm_1 | ln_1_land_226_lpi_1_dfm_1 | ln_1_land_227_lpi_1_dfm_1
          | ln_1_land_229_lpi_1_dfm_1 | ln_1_land_230_lpi_1_dfm_1 | ln_1_land_232_lpi_1_dfm_1
          | ln_1_land_233_lpi_1_dfm_1 | ln_1_land_239_lpi_1_dfm_1 | ln_1_land_240_lpi_1_dfm_1
          | ln_1_land_242_lpi_1_dfm_1 | ln_1_land_244_lpi_1_dfm_1;
      ln_1_ln_1_mux1h_118_psp_1_2 <= (((~((~((((~(((~(ln_1_nor_5_cse_1 | ln_1_and_2_ssc_1
          | ln_1_land_6_lpi_1_dfm_1)) & (~(ln_1_and_4_ssc_1 | ln_1_land_8_lpi_1_dfm_1
          | ln_1_land_10_lpi_1_dfm_1 | ln_1_land_12_lpi_1_dfm_1 | ln_1_land_13_lpi_1_dfm_1
          | ln_1_land_15_lpi_1_dfm_1 | ln_1_land_18_lpi_1_dfm_1 | ln_1_land_19_lpi_1_dfm_1
          | ln_1_land_21_lpi_1_dfm_1 | ln_1_land_22_lpi_1_dfm_1 | ln_1_land_25_lpi_1_dfm_1
          | ln_1_land_26_lpi_1_dfm_1 | ln_1_land_30_lpi_1_dfm_1 | ln_1_land_31_lpi_1_dfm_1
          | ln_1_land_32_lpi_1_dfm_1 | ln_1_land_38_lpi_1_dfm_1 | ln_1_land_39_lpi_1_dfm_1
          | ln_1_land_40_lpi_1_dfm_1 | ln_1_land_41_lpi_1_dfm_1 | ln_1_land_42_lpi_1_dfm_1
          | ln_1_land_43_lpi_1_dfm_1 | ln_1_land_44_lpi_1_dfm_1 | ln_1_land_45_lpi_1_dfm_1
          | ln_1_land_46_lpi_1_dfm_1))) | ln_1_land_9_lpi_1_dfm_1 | ln_1_land_11_lpi_1_dfm_1
          | ln_1_land_14_lpi_1_dfm_1 | ln_1_land_16_lpi_1_dfm_1 | ln_1_land_17_lpi_1_dfm_1
          | ln_1_land_20_lpi_1_dfm_1 | ln_1_land_23_lpi_1_dfm_1 | ln_1_land_24_lpi_1_dfm_1
          | ln_1_land_27_lpi_1_dfm_1 | ln_1_land_28_lpi_1_dfm_1 | ln_1_land_29_lpi_1_dfm_1
          | ln_1_land_33_lpi_1_dfm_1 | ln_1_land_34_lpi_1_dfm_1 | ln_1_land_35_lpi_1_dfm_1
          | ln_1_land_36_lpi_1_dfm_1 | ln_1_land_37_lpi_1_dfm_1 | ln_1_land_47_lpi_1_dfm_1
          | ln_1_land_48_lpi_1_dfm_1 | ln_1_land_49_lpi_1_dfm_1 | ln_1_if_50_ln_1_if_50_and_seb_1))
          | ln_1_land_51_lpi_1_dfm_1 | ln_1_land_52_lpi_1_dfm_1) & (~(ln_1_land_54_lpi_1_dfm_1
          | ln_1_land_55_lpi_1_dfm_1 | ln_1_land_58_lpi_1_dfm_1 | ln_1_land_59_lpi_1_dfm_1
          | ln_1_land_61_lpi_1_dfm_1 | ln_1_land_62_lpi_1_dfm_1 | ln_1_land_64_lpi_1_dfm_1
          | ln_1_land_66_lpi_1_dfm_1 | ln_1_land_68_lpi_1_dfm_1 | ln_1_land_70_lpi_1_dfm_1
          | ln_1_land_72_lpi_1_dfm_1 | ln_1_land_75_lpi_1_dfm_1 | ln_1_land_78_lpi_1_dfm_1
          | ln_1_land_79_lpi_1_dfm_1 | ln_1_land_80_lpi_1_dfm_1 | ln_1_land_89_lpi_1_dfm_1
          | ln_1_land_90_lpi_1_dfm_1 | ln_1_land_93_lpi_1_dfm_1 | ln_1_land_94_lpi_1_dfm_1
          | ln_1_land_96_lpi_1_dfm_1 | ln_1_land_98_lpi_1_dfm_1 | ln_1_land_101_lpi_1_dfm_1
          | ln_1_land_106_lpi_1_dfm_1 | ln_1_land_110_lpi_1_dfm_1 | ln_1_land_111_lpi_1_dfm_1
          | ln_1_land_113_lpi_1_dfm_1 | ln_1_land_115_lpi_1_dfm_1 | ln_1_land_116_lpi_1_dfm_1
          | ln_1_land_120_lpi_1_dfm_1 | ln_1_land_123_lpi_1_dfm_1 | ln_1_land_125_lpi_1_dfm_1
          | ln_1_land_126_lpi_1_dfm_1 | ln_1_land_129_lpi_1_dfm_1 | ln_1_land_132_lpi_1_dfm_1
          | ln_1_land_133_lpi_1_dfm_1 | ln_1_land_136_lpi_1_dfm_1 | ln_1_land_137_lpi_1_dfm_1
          | ln_1_land_138_lpi_1_dfm_1))) | ln_1_and_48_ssc_1 | ln_1_land_56_lpi_1_dfm_1
          | ln_1_land_57_lpi_1_dfm_1 | ln_1_land_60_lpi_1_dfm_1 | ln_1_land_63_lpi_1_dfm_1
          | ln_1_land_65_lpi_1_dfm_1 | ln_1_land_67_lpi_1_dfm_1 | ln_1_land_69_lpi_1_dfm_1
          | ln_1_land_71_lpi_1_dfm_1 | ln_1_land_73_lpi_1_dfm_1 | ln_1_land_74_lpi_1_dfm_1
          | ln_1_land_76_lpi_1_dfm_1 | ln_1_land_77_lpi_1_dfm_1 | ln_1_land_81_lpi_1_dfm_1
          | ln_1_land_82_lpi_1_dfm_1 | ln_1_land_83_lpi_1_dfm_1 | ln_1_land_84_lpi_1_dfm_1
          | ln_1_land_85_lpi_1_dfm_1 | ln_1_land_86_lpi_1_dfm_1 | ln_1_land_87_lpi_1_dfm_1
          | ln_1_land_88_lpi_1_dfm_1 | ln_1_land_91_lpi_1_dfm_1 | ln_1_land_92_lpi_1_dfm_1
          | ln_1_land_95_lpi_1_dfm_1 | ln_1_land_97_lpi_1_dfm_1 | ln_1_land_99_lpi_1_dfm_1
          | ln_1_land_100_lpi_1_dfm_1 | ln_1_land_102_lpi_1_dfm_1 | ln_1_land_103_lpi_1_dfm_1
          | ln_1_land_104_lpi_1_dfm_1 | ln_1_land_105_lpi_1_dfm_1 | ln_1_land_107_lpi_1_dfm_1
          | ln_1_land_108_lpi_1_dfm_1 | ln_1_land_109_lpi_1_dfm_1 | ln_1_land_112_lpi_1_dfm_1
          | ln_1_land_114_lpi_1_dfm_1 | ln_1_land_117_lpi_1_dfm_1 | ln_1_land_118_lpi_1_dfm_1
          | ln_1_land_119_lpi_1_dfm_1 | ln_1_land_121_lpi_1_dfm_1 | ln_1_land_122_lpi_1_dfm_1
          | ln_1_land_124_lpi_1_dfm_1 | ln_1_land_127_lpi_1_dfm_1 | ln_1_land_128_lpi_1_dfm_1
          | ln_1_land_130_lpi_1_dfm_1 | ln_1_land_131_lpi_1_dfm_1 | ln_1_land_134_lpi_1_dfm_1
          | ln_1_land_135_lpi_1_dfm_1 | ln_1_land_139_lpi_1_dfm_1 | ln_1_land_140_lpi_1_dfm_1))
          | ln_1_land_142_lpi_1_dfm_1)) | ln_1_land_141_lpi_1_dfm_1) & ln_1_nor_3_cse_1
          & (~(ln_1_and_140_ssc_1 | ln_1_land_146_lpi_1_dfm_1 | ln_1_land_156_lpi_1_dfm_1
          | ln_1_land_157_lpi_1_dfm_1 | ln_1_land_158_lpi_1_dfm_1 | ln_1_land_159_lpi_1_dfm_1
          | ln_1_land_163_lpi_1_dfm_1 | ln_1_land_164_lpi_1_dfm_1 | ln_1_land_165_lpi_1_dfm_1
          | ln_1_land_167_lpi_1_dfm_1 | ln_1_land_168_lpi_1_dfm_1 | ln_1_land_171_lpi_1_dfm_1
          | ln_1_land_173_lpi_1_dfm_1 | ln_1_land_176_lpi_1_dfm_1 | ln_1_land_178_lpi_1_dfm_1
          | ln_1_land_179_lpi_1_dfm_1 | ln_1_land_181_lpi_1_dfm_1 | ln_1_land_183_lpi_1_dfm_1
          | ln_1_land_184_lpi_1_dfm_1 | ln_1_land_187_lpi_1_dfm_1 | ln_1_land_188_lpi_1_dfm_1
          | ln_1_land_189_lpi_1_dfm_1 | ln_1_land_199_lpi_1_dfm_1 | ln_1_land_200_lpi_1_dfm_1
          | ln_1_land_203_lpi_1_dfm_1 | ln_1_land_205_lpi_1_dfm_1 | ln_1_land_207_lpi_1_dfm_1
          | ln_1_land_209_lpi_1_dfm_1 | ln_1_land_210_lpi_1_dfm_1 | ln_1_land_213_lpi_1_dfm_1
          | ln_1_land_214_lpi_1_dfm_1 | ln_1_land_215_lpi_1_dfm_1 | ln_1_land_216_lpi_1_dfm_1
          | ln_1_land_217_lpi_1_dfm_1 | ln_1_land_220_lpi_1_dfm_1 | ln_1_land_221_lpi_1_dfm_1
          | ln_1_land_223_lpi_1_dfm_1 | ln_1_land_224_lpi_1_dfm_1 | ln_1_land_227_lpi_1_dfm_1
          | ln_1_land_228_lpi_1_dfm_1 | ln_1_land_229_lpi_1_dfm_1 | ln_1_land_232_lpi_1_dfm_1
          | ln_1_land_234_lpi_1_dfm_1 | ln_1_land_235_lpi_1_dfm_1 | ln_1_land_236_lpi_1_dfm_1
          | ln_1_land_237_lpi_1_dfm_1 | ln_1_land_238_lpi_1_dfm_1 | ln_1_land_240_lpi_1_dfm_1)))
          | ln_1_land_147_lpi_1_dfm_1 | ln_1_land_148_lpi_1_dfm_1 | ln_1_land_149_lpi_1_dfm_1
          | ln_1_land_150_lpi_1_dfm_1 | ln_1_land_151_lpi_1_dfm_1 | ln_1_land_152_lpi_1_dfm_1
          | ln_1_land_153_lpi_1_dfm_1 | ln_1_land_154_lpi_1_dfm_1 | ln_1_land_155_lpi_1_dfm_1
          | ln_1_land_160_lpi_1_dfm_1 | ln_1_land_161_lpi_1_dfm_1 | ln_1_land_162_lpi_1_dfm_1
          | ln_1_land_166_lpi_1_dfm_1 | ln_1_land_169_lpi_1_dfm_1 | ln_1_land_170_lpi_1_dfm_1
          | ln_1_land_172_lpi_1_dfm_1 | ln_1_land_174_lpi_1_dfm_1 | ln_1_land_175_lpi_1_dfm_1
          | ln_1_land_177_lpi_1_dfm_1 | ln_1_land_180_lpi_1_dfm_1 | ln_1_land_182_lpi_1_dfm_1
          | ln_1_land_185_lpi_1_dfm_1 | ln_1_land_186_lpi_1_dfm_1 | ln_1_land_190_lpi_1_dfm_1
          | ln_1_land_191_lpi_1_dfm_1 | ln_1_land_192_lpi_1_dfm_1 | ln_1_land_193_lpi_1_dfm_1
          | ln_1_land_194_lpi_1_dfm_1 | ln_1_land_195_lpi_1_dfm_1 | ln_1_land_196_lpi_1_dfm_1
          | ln_1_land_197_lpi_1_dfm_1 | ln_1_land_198_lpi_1_dfm_1 | ln_1_land_201_lpi_1_dfm_1
          | ln_1_land_202_lpi_1_dfm_1 | ln_1_land_204_lpi_1_dfm_1 | ln_1_land_206_lpi_1_dfm_1
          | ln_1_land_208_lpi_1_dfm_1 | ln_1_land_211_lpi_1_dfm_1 | ln_1_land_212_lpi_1_dfm_1
          | ln_1_land_218_lpi_1_dfm_1 | ln_1_land_219_lpi_1_dfm_1 | ln_1_land_222_lpi_1_dfm_1
          | ln_1_land_225_lpi_1_dfm_1 | ln_1_land_226_lpi_1_dfm_1 | ln_1_land_230_lpi_1_dfm_1
          | ln_1_land_231_lpi_1_dfm_1 | ln_1_land_233_lpi_1_dfm_1 | ln_1_land_239_lpi_1_dfm_1
          | ln_1_land_241_lpi_1_dfm_1 | ln_1_land_242_lpi_1_dfm_1 | ln_1_land_243_lpi_1_dfm_1
          | ln_1_land_244_lpi_1_dfm_1;
      ln_1_ln_1_mux1h_118_psp_1_1 <= (((~((~((~((~((((~(((ln_1_land_4_lpi_1_dfm_1
          | ln_1_and_2_ssc_1 | ln_1_land_6_lpi_1_dfm_1) & (~(ln_1_land_8_lpi_1_dfm_1
          | ln_1_land_9_lpi_1_dfm_1 | ln_1_land_10_lpi_1_dfm_1 | ln_1_land_13_lpi_1_dfm_1
          | ln_1_land_14_lpi_1_dfm_1 | ln_1_land_17_lpi_1_dfm_1 | ln_1_land_19_lpi_1_dfm_1
          | ln_1_land_20_lpi_1_dfm_1 | ln_1_land_22_lpi_1_dfm_1 | ln_1_land_24_lpi_1_dfm_1
          | ln_1_land_26_lpi_1_dfm_1 | ln_1_land_29_lpi_1_dfm_1 | ln_1_land_31_lpi_1_dfm_1
          | ln_1_land_32_lpi_1_dfm_1 | ln_1_land_35_lpi_1_dfm_1 | ln_1_land_36_lpi_1_dfm_1
          | ln_1_land_37_lpi_1_dfm_1 | ln_1_land_47_lpi_1_dfm_1 | ln_1_land_48_lpi_1_dfm_1)))
          | ln_1_and_4_ssc_1 | ln_1_land_11_lpi_1_dfm_1 | ln_1_land_12_lpi_1_dfm_1
          | ln_1_land_15_lpi_1_dfm_1 | ln_1_land_16_lpi_1_dfm_1 | ln_1_land_18_lpi_1_dfm_1
          | ln_1_land_21_lpi_1_dfm_1 | ln_1_land_23_lpi_1_dfm_1 | ln_1_land_25_lpi_1_dfm_1
          | ln_1_land_27_lpi_1_dfm_1 | ln_1_land_28_lpi_1_dfm_1 | ln_1_land_30_lpi_1_dfm_1
          | ln_1_land_33_lpi_1_dfm_1 | ln_1_land_34_lpi_1_dfm_1 | ln_1_land_38_lpi_1_dfm_1
          | ln_1_land_39_lpi_1_dfm_1 | ln_1_land_40_lpi_1_dfm_1 | ln_1_land_41_lpi_1_dfm_1
          | ln_1_land_42_lpi_1_dfm_1 | ln_1_land_43_lpi_1_dfm_1 | ln_1_land_44_lpi_1_dfm_1
          | ln_1_land_45_lpi_1_dfm_1 | ln_1_land_46_lpi_1_dfm_1 | ln_1_land_49_lpi_1_dfm_1
          | ln_1_if_50_ln_1_if_50_and_seb_1)) | ln_1_land_51_lpi_1_dfm_1 | ln_1_land_52_lpi_1_dfm_1)
          & (~(ln_1_and_48_ssc_1 | ln_1_land_55_lpi_1_dfm_1 | ln_1_land_57_lpi_1_dfm_1
          | ln_1_land_59_lpi_1_dfm_1 | ln_1_land_62_lpi_1_dfm_1 | ln_1_land_63_lpi_1_dfm_1
          | ln_1_land_72_lpi_1_dfm_1 | ln_1_land_73_lpi_1_dfm_1 | ln_1_land_75_lpi_1_dfm_1
          | ln_1_land_76_lpi_1_dfm_1 | ln_1_land_78_lpi_1_dfm_1 | ln_1_land_79_lpi_1_dfm_1
          | ln_1_land_81_lpi_1_dfm_1 | ln_1_land_82_lpi_1_dfm_1 | ln_1_land_83_lpi_1_dfm_1
          | ln_1_land_84_lpi_1_dfm_1 | ln_1_land_85_lpi_1_dfm_1 | ln_1_land_86_lpi_1_dfm_1
          | ln_1_land_87_lpi_1_dfm_1 | ln_1_land_88_lpi_1_dfm_1 | ln_1_land_90_lpi_1_dfm_1
          | ln_1_land_92_lpi_1_dfm_1 | ln_1_land_94_lpi_1_dfm_1 | ln_1_land_95_lpi_1_dfm_1
          | ln_1_land_96_lpi_1_dfm_1 | ln_1_land_97_lpi_1_dfm_1 | ln_1_land_98_lpi_1_dfm_1
          | ln_1_land_99_lpi_1_dfm_1 | ln_1_land_102_lpi_1_dfm_1 | ln_1_land_106_lpi_1_dfm_1
          | ln_1_land_109_lpi_1_dfm_1 | ln_1_land_111_lpi_1_dfm_1 | ln_1_land_115_lpi_1_dfm_1
          | ln_1_land_117_lpi_1_dfm_1 | ln_1_land_120_lpi_1_dfm_1 | ln_1_land_121_lpi_1_dfm_1
          | ln_1_land_124_lpi_1_dfm_1 | ln_1_land_125_lpi_1_dfm_1 | ln_1_land_127_lpi_1_dfm_1
          | ln_1_land_130_lpi_1_dfm_1 | ln_1_land_132_lpi_1_dfm_1 | ln_1_land_134_lpi_1_dfm_1
          | ln_1_land_136_lpi_1_dfm_1 | ln_1_land_137_lpi_1_dfm_1 | ln_1_land_139_lpi_1_dfm_1)))
          | ln_1_land_54_lpi_1_dfm_1 | ln_1_land_56_lpi_1_dfm_1 | ln_1_land_58_lpi_1_dfm_1
          | ln_1_land_60_lpi_1_dfm_1 | ln_1_land_61_lpi_1_dfm_1 | ln_1_land_64_lpi_1_dfm_1
          | ln_1_land_65_lpi_1_dfm_1 | ln_1_land_66_lpi_1_dfm_1 | ln_1_land_67_lpi_1_dfm_1
          | ln_1_land_68_lpi_1_dfm_1 | ln_1_land_69_lpi_1_dfm_1 | ln_1_land_70_lpi_1_dfm_1
          | ln_1_land_71_lpi_1_dfm_1 | ln_1_land_74_lpi_1_dfm_1 | ln_1_land_77_lpi_1_dfm_1
          | ln_1_land_80_lpi_1_dfm_1 | ln_1_land_89_lpi_1_dfm_1 | ln_1_land_91_lpi_1_dfm_1
          | ln_1_land_93_lpi_1_dfm_1 | ln_1_land_100_lpi_1_dfm_1 | ln_1_land_101_lpi_1_dfm_1
          | ln_1_land_103_lpi_1_dfm_1 | ln_1_land_104_lpi_1_dfm_1 | ln_1_land_105_lpi_1_dfm_1
          | ln_1_land_107_lpi_1_dfm_1 | ln_1_land_108_lpi_1_dfm_1 | ln_1_land_110_lpi_1_dfm_1
          | ln_1_land_112_lpi_1_dfm_1 | ln_1_land_113_lpi_1_dfm_1 | ln_1_land_114_lpi_1_dfm_1
          | ln_1_land_116_lpi_1_dfm_1 | ln_1_land_118_lpi_1_dfm_1 | ln_1_land_119_lpi_1_dfm_1
          | ln_1_land_122_lpi_1_dfm_1 | ln_1_land_123_lpi_1_dfm_1 | ln_1_land_126_lpi_1_dfm_1
          | ln_1_land_128_lpi_1_dfm_1 | ln_1_land_129_lpi_1_dfm_1 | ln_1_land_131_lpi_1_dfm_1
          | ln_1_land_133_lpi_1_dfm_1 | ln_1_land_135_lpi_1_dfm_1 | ln_1_land_138_lpi_1_dfm_1
          | ln_1_land_140_lpi_1_dfm_1)) | ln_1_land_142_lpi_1_dfm_1)) | ln_1_land_141_lpi_1_dfm_1))
          | ln_1_and_138_ssc_1)) | ln_1_land_144_lpi_1_dfm_1) & (~(ln_1_land_147_lpi_1_dfm_1
          | ln_1_land_148_lpi_1_dfm_1 | ln_1_land_149_lpi_1_dfm_1 | ln_1_land_150_lpi_1_dfm_1
          | ln_1_land_151_lpi_1_dfm_1 | ln_1_land_152_lpi_1_dfm_1 | ln_1_land_153_lpi_1_dfm_1
          | ln_1_land_154_lpi_1_dfm_1 | ln_1_land_155_lpi_1_dfm_1 | ln_1_land_159_lpi_1_dfm_1
          | ln_1_land_162_lpi_1_dfm_1 | ln_1_land_164_lpi_1_dfm_1 | ln_1_land_165_lpi_1_dfm_1
          | ln_1_land_168_lpi_1_dfm_1 | ln_1_land_170_lpi_1_dfm_1 | ln_1_land_171_lpi_1_dfm_1
          | ln_1_land_175_lpi_1_dfm_1 | ln_1_land_176_lpi_1_dfm_1 | ln_1_land_177_lpi_1_dfm_1
          | ln_1_land_178_lpi_1_dfm_1 | ln_1_land_182_lpi_1_dfm_1 | ln_1_land_183_lpi_1_dfm_1
          | ln_1_land_185_lpi_1_dfm_1 | ln_1_land_187_lpi_1_dfm_1 | ln_1_land_190_lpi_1_dfm_1
          | ln_1_land_191_lpi_1_dfm_1 | ln_1_land_197_lpi_1_dfm_1 | ln_1_land_198_lpi_1_dfm_1
          | ln_1_land_200_lpi_1_dfm_1 | ln_1_land_202_lpi_1_dfm_1 | ln_1_land_203_lpi_1_dfm_1
          | ln_1_land_209_lpi_1_dfm_1 | ln_1_land_211_lpi_1_dfm_1 | ln_1_land_213_lpi_1_dfm_1
          | ln_1_land_214_lpi_1_dfm_1 | ln_1_land_215_lpi_1_dfm_1 | ln_1_land_216_lpi_1_dfm_1
          | ln_1_land_217_lpi_1_dfm_1 | ln_1_land_219_lpi_1_dfm_1 | ln_1_land_221_lpi_1_dfm_1
          | ln_1_land_222_lpi_1_dfm_1 | ln_1_land_223_lpi_1_dfm_1 | ln_1_land_225_lpi_1_dfm_1
          | ln_1_land_227_lpi_1_dfm_1 | ln_1_land_228_lpi_1_dfm_1 | ln_1_land_229_lpi_1_dfm_1
          | ln_1_land_231_lpi_1_dfm_1 | ln_1_land_232_lpi_1_dfm_1 | ln_1_land_233_lpi_1_dfm_1
          | ln_1_land_234_lpi_1_dfm_1 | ln_1_land_238_lpi_1_dfm_1 | ln_1_land_244_lpi_1_dfm_1)))
          | ln_1_and_140_ssc_1 | ln_1_land_146_lpi_1_dfm_1 | ln_1_land_156_lpi_1_dfm_1
          | ln_1_land_157_lpi_1_dfm_1 | ln_1_land_158_lpi_1_dfm_1 | ln_1_land_160_lpi_1_dfm_1
          | ln_1_land_161_lpi_1_dfm_1 | ln_1_land_163_lpi_1_dfm_1 | ln_1_land_166_lpi_1_dfm_1
          | ln_1_land_167_lpi_1_dfm_1 | ln_1_land_169_lpi_1_dfm_1 | ln_1_land_172_lpi_1_dfm_1
          | ln_1_land_173_lpi_1_dfm_1 | ln_1_land_174_lpi_1_dfm_1 | ln_1_land_179_lpi_1_dfm_1
          | ln_1_land_180_lpi_1_dfm_1 | ln_1_land_181_lpi_1_dfm_1 | ln_1_land_184_lpi_1_dfm_1
          | ln_1_land_186_lpi_1_dfm_1 | ln_1_land_188_lpi_1_dfm_1 | ln_1_land_189_lpi_1_dfm_1
          | ln_1_land_192_lpi_1_dfm_1 | ln_1_land_193_lpi_1_dfm_1 | ln_1_land_194_lpi_1_dfm_1
          | ln_1_land_195_lpi_1_dfm_1 | ln_1_land_196_lpi_1_dfm_1 | ln_1_land_199_lpi_1_dfm_1
          | ln_1_land_201_lpi_1_dfm_1 | ln_1_land_204_lpi_1_dfm_1 | ln_1_land_205_lpi_1_dfm_1
          | ln_1_land_206_lpi_1_dfm_1 | ln_1_land_207_lpi_1_dfm_1 | ln_1_land_208_lpi_1_dfm_1
          | ln_1_land_210_lpi_1_dfm_1 | ln_1_land_212_lpi_1_dfm_1 | ln_1_land_218_lpi_1_dfm_1
          | ln_1_land_220_lpi_1_dfm_1 | ln_1_land_224_lpi_1_dfm_1 | ln_1_land_226_lpi_1_dfm_1
          | ln_1_land_230_lpi_1_dfm_1 | ln_1_land_235_lpi_1_dfm_1 | ln_1_land_236_lpi_1_dfm_1
          | ln_1_land_237_lpi_1_dfm_1 | ln_1_land_239_lpi_1_dfm_1 | ln_1_land_240_lpi_1_dfm_1
          | ln_1_land_241_lpi_1_dfm_1 | ln_1_land_242_lpi_1_dfm_1 | ln_1_land_243_lpi_1_dfm_1;
      ln_1_ln_1_mux1h_118_psp_1_0 <= (((~((~((~((~((((~((ln_1_nor_1_cse_1 & (~(ln_1_land_8_lpi_1_dfm_1
          | ln_1_land_9_lpi_1_dfm_1 | ln_1_land_11_lpi_1_dfm_1 | ln_1_land_13_lpi_1_dfm_1
          | ln_1_land_15_lpi_1_dfm_1 | ln_1_land_18_lpi_1_dfm_1 | ln_1_land_19_lpi_1_dfm_1
          | ln_1_land_28_lpi_1_dfm_1 | ln_1_land_29_lpi_1_dfm_1 | ln_1_land_32_lpi_1_dfm_1
          | ln_1_land_34_lpi_1_dfm_1 | ln_1_land_37_lpi_1_dfm_1 | ln_1_land_41_lpi_1_dfm_1
          | ln_1_land_42_lpi_1_dfm_1 | ln_1_land_43_lpi_1_dfm_1 | ln_1_land_47_lpi_1_dfm_1
          | ln_1_land_49_lpi_1_dfm_1))) | ln_1_and_4_ssc_1 | ln_1_land_10_lpi_1_dfm_1
          | ln_1_land_12_lpi_1_dfm_1 | ln_1_land_14_lpi_1_dfm_1 | ln_1_land_16_lpi_1_dfm_1
          | ln_1_land_17_lpi_1_dfm_1 | ln_1_land_20_lpi_1_dfm_1 | ln_1_land_21_lpi_1_dfm_1
          | ln_1_land_22_lpi_1_dfm_1 | ln_1_land_23_lpi_1_dfm_1 | ln_1_land_24_lpi_1_dfm_1
          | ln_1_land_25_lpi_1_dfm_1 | ln_1_land_26_lpi_1_dfm_1 | ln_1_land_27_lpi_1_dfm_1
          | ln_1_land_30_lpi_1_dfm_1 | ln_1_land_31_lpi_1_dfm_1 | ln_1_land_33_lpi_1_dfm_1
          | ln_1_land_35_lpi_1_dfm_1 | ln_1_land_36_lpi_1_dfm_1 | ln_1_land_38_lpi_1_dfm_1
          | ln_1_land_39_lpi_1_dfm_1 | ln_1_land_40_lpi_1_dfm_1 | ln_1_land_44_lpi_1_dfm_1
          | ln_1_land_45_lpi_1_dfm_1 | ln_1_land_46_lpi_1_dfm_1 | ln_1_land_48_lpi_1_dfm_1
          | ln_1_if_50_ln_1_if_50_and_seb_1 | ln_1_land_52_lpi_1_dfm_1)) | ln_1_land_51_lpi_1_dfm_1)
          & (~(ln_1_and_48_ssc_1 | ln_1_land_60_lpi_1_dfm_1 | ln_1_land_62_lpi_1_dfm_1
          | ln_1_land_64_lpi_1_dfm_1 | ln_1_land_71_lpi_1_dfm_1 | ln_1_land_73_lpi_1_dfm_1
          | ln_1_land_76_lpi_1_dfm_1 | ln_1_land_77_lpi_1_dfm_1 | ln_1_land_78_lpi_1_dfm_1
          | ln_1_land_81_lpi_1_dfm_1 | ln_1_land_88_lpi_1_dfm_1 | ln_1_land_94_lpi_1_dfm_1
          | ln_1_land_99_lpi_1_dfm_1 | ln_1_land_101_lpi_1_dfm_1 | ln_1_land_102_lpi_1_dfm_1
          | ln_1_land_103_lpi_1_dfm_1 | ln_1_land_106_lpi_1_dfm_1 | ln_1_land_108_lpi_1_dfm_1
          | ln_1_land_112_lpi_1_dfm_1 | ln_1_land_113_lpi_1_dfm_1 | ln_1_land_114_lpi_1_dfm_1
          | ln_1_land_118_lpi_1_dfm_1 | ln_1_land_119_lpi_1_dfm_1 | ln_1_land_121_lpi_1_dfm_1
          | ln_1_land_123_lpi_1_dfm_1 | ln_1_land_125_lpi_1_dfm_1 | ln_1_land_126_lpi_1_dfm_1
          | ln_1_land_129_lpi_1_dfm_1 | ln_1_land_130_lpi_1_dfm_1 | ln_1_land_131_lpi_1_dfm_1
          | ln_1_land_132_lpi_1_dfm_1 | ln_1_land_133_lpi_1_dfm_1 | ln_1_land_134_lpi_1_dfm_1
          | ln_1_land_135_lpi_1_dfm_1 | ln_1_land_136_lpi_1_dfm_1 | ln_1_land_139_lpi_1_dfm_1
          | ln_1_land_140_lpi_1_dfm_1))) | ln_1_land_54_lpi_1_dfm_1 | ln_1_land_55_lpi_1_dfm_1
          | ln_1_land_56_lpi_1_dfm_1 | ln_1_land_57_lpi_1_dfm_1 | ln_1_land_58_lpi_1_dfm_1
          | ln_1_land_59_lpi_1_dfm_1 | ln_1_land_61_lpi_1_dfm_1 | ln_1_land_63_lpi_1_dfm_1
          | ln_1_land_65_lpi_1_dfm_1 | ln_1_land_66_lpi_1_dfm_1 | ln_1_land_67_lpi_1_dfm_1
          | ln_1_land_68_lpi_1_dfm_1 | ln_1_land_69_lpi_1_dfm_1 | ln_1_land_70_lpi_1_dfm_1
          | ln_1_land_72_lpi_1_dfm_1 | ln_1_land_74_lpi_1_dfm_1 | ln_1_land_75_lpi_1_dfm_1
          | ln_1_land_79_lpi_1_dfm_1 | ln_1_land_80_lpi_1_dfm_1 | ln_1_land_82_lpi_1_dfm_1
          | ln_1_land_83_lpi_1_dfm_1 | ln_1_land_84_lpi_1_dfm_1 | ln_1_land_85_lpi_1_dfm_1
          | ln_1_land_86_lpi_1_dfm_1 | ln_1_land_87_lpi_1_dfm_1 | ln_1_land_89_lpi_1_dfm_1
          | ln_1_land_90_lpi_1_dfm_1 | ln_1_land_91_lpi_1_dfm_1 | ln_1_land_92_lpi_1_dfm_1
          | ln_1_land_93_lpi_1_dfm_1 | ln_1_land_95_lpi_1_dfm_1 | ln_1_land_96_lpi_1_dfm_1
          | ln_1_land_97_lpi_1_dfm_1 | ln_1_land_98_lpi_1_dfm_1 | ln_1_land_100_lpi_1_dfm_1
          | ln_1_land_104_lpi_1_dfm_1 | ln_1_land_105_lpi_1_dfm_1 | ln_1_land_107_lpi_1_dfm_1
          | ln_1_land_109_lpi_1_dfm_1 | ln_1_land_110_lpi_1_dfm_1 | ln_1_land_111_lpi_1_dfm_1
          | ln_1_land_115_lpi_1_dfm_1 | ln_1_land_116_lpi_1_dfm_1 | ln_1_land_117_lpi_1_dfm_1
          | ln_1_land_120_lpi_1_dfm_1 | ln_1_land_122_lpi_1_dfm_1 | ln_1_land_124_lpi_1_dfm_1
          | ln_1_land_127_lpi_1_dfm_1 | ln_1_land_128_lpi_1_dfm_1 | ln_1_land_137_lpi_1_dfm_1
          | ln_1_land_138_lpi_1_dfm_1)) | ln_1_land_142_lpi_1_dfm_1)) | ln_1_land_141_lpi_1_dfm_1))
          | ln_1_land_144_lpi_1_dfm_1)) | ln_1_and_138_ssc_1) & (~(ln_1_land_147_lpi_1_dfm_1
          | ln_1_land_148_lpi_1_dfm_1 | ln_1_land_154_lpi_1_dfm_1 | ln_1_land_155_lpi_1_dfm_1
          | ln_1_land_157_lpi_1_dfm_1 | ln_1_land_158_lpi_1_dfm_1 | ln_1_land_161_lpi_1_dfm_1
          | ln_1_land_165_lpi_1_dfm_1 | ln_1_land_166_lpi_1_dfm_1 | ln_1_land_169_lpi_1_dfm_1
          | ln_1_land_170_lpi_1_dfm_1 | ln_1_land_172_lpi_1_dfm_1 | ln_1_land_175_lpi_1_dfm_1
          | ln_1_land_176_lpi_1_dfm_1 | ln_1_land_177_lpi_1_dfm_1 | ln_1_land_178_lpi_1_dfm_1
          | ln_1_land_181_lpi_1_dfm_1 | ln_1_land_183_lpi_1_dfm_1 | ln_1_land_184_lpi_1_dfm_1
          | ln_1_land_187_lpi_1_dfm_1 | ln_1_land_188_lpi_1_dfm_1 | ln_1_land_192_lpi_1_dfm_1
          | ln_1_land_193_lpi_1_dfm_1 | ln_1_land_194_lpi_1_dfm_1 | ln_1_land_195_lpi_1_dfm_1
          | ln_1_land_196_lpi_1_dfm_1 | ln_1_land_198_lpi_1_dfm_1 | ln_1_land_199_lpi_1_dfm_1
          | ln_1_land_200_lpi_1_dfm_1 | ln_1_land_201_lpi_1_dfm_1 | ln_1_land_202_lpi_1_dfm_1
          | ln_1_land_204_lpi_1_dfm_1 | ln_1_land_207_lpi_1_dfm_1 | ln_1_land_208_lpi_1_dfm_1
          | ln_1_land_213_lpi_1_dfm_1 | ln_1_land_217_lpi_1_dfm_1 | ln_1_land_221_lpi_1_dfm_1
          | ln_1_land_222_lpi_1_dfm_1 | ln_1_land_223_lpi_1_dfm_1 | ln_1_land_227_lpi_1_dfm_1
          | ln_1_land_228_lpi_1_dfm_1 | ln_1_land_229_lpi_1_dfm_1 | ln_1_land_230_lpi_1_dfm_1
          | ln_1_land_231_lpi_1_dfm_1 | ln_1_land_234_lpi_1_dfm_1 | ln_1_land_235_lpi_1_dfm_1
          | ln_1_land_241_lpi_1_dfm_1))) | ln_1_and_140_ssc_1 | ln_1_land_146_lpi_1_dfm_1
          | ln_1_land_149_lpi_1_dfm_1 | ln_1_land_150_lpi_1_dfm_1 | ln_1_land_151_lpi_1_dfm_1
          | ln_1_land_152_lpi_1_dfm_1 | ln_1_land_153_lpi_1_dfm_1 | ln_1_land_156_lpi_1_dfm_1
          | ln_1_land_159_lpi_1_dfm_1 | ln_1_land_160_lpi_1_dfm_1 | ln_1_land_162_lpi_1_dfm_1
          | ln_1_land_163_lpi_1_dfm_1 | ln_1_land_164_lpi_1_dfm_1 | ln_1_land_167_lpi_1_dfm_1
          | ln_1_land_168_lpi_1_dfm_1 | ln_1_land_171_lpi_1_dfm_1 | ln_1_land_173_lpi_1_dfm_1
          | ln_1_land_174_lpi_1_dfm_1 | ln_1_land_179_lpi_1_dfm_1 | ln_1_land_180_lpi_1_dfm_1
          | ln_1_land_182_lpi_1_dfm_1 | ln_1_land_185_lpi_1_dfm_1 | ln_1_land_186_lpi_1_dfm_1
          | ln_1_land_189_lpi_1_dfm_1 | ln_1_land_190_lpi_1_dfm_1 | ln_1_land_191_lpi_1_dfm_1
          | ln_1_land_197_lpi_1_dfm_1 | ln_1_land_203_lpi_1_dfm_1 | ln_1_land_205_lpi_1_dfm_1
          | ln_1_land_206_lpi_1_dfm_1 | ln_1_land_209_lpi_1_dfm_1 | ln_1_land_210_lpi_1_dfm_1
          | ln_1_land_211_lpi_1_dfm_1 | ln_1_land_212_lpi_1_dfm_1 | ln_1_land_214_lpi_1_dfm_1
          | ln_1_land_215_lpi_1_dfm_1 | ln_1_land_216_lpi_1_dfm_1 | ln_1_land_218_lpi_1_dfm_1
          | ln_1_land_219_lpi_1_dfm_1 | ln_1_land_220_lpi_1_dfm_1 | ln_1_land_224_lpi_1_dfm_1
          | ln_1_land_225_lpi_1_dfm_1 | ln_1_land_226_lpi_1_dfm_1 | ln_1_land_232_lpi_1_dfm_1
          | ln_1_land_233_lpi_1_dfm_1 | ln_1_land_236_lpi_1_dfm_1 | ln_1_land_237_lpi_1_dfm_1
          | ln_1_land_238_lpi_1_dfm_1 | ln_1_land_239_lpi_1_dfm_1 | ln_1_land_240_lpi_1_dfm_1
          | ln_1_land_242_lpi_1_dfm_1 | ln_1_land_243_lpi_1_dfm_1 | ln_1_land_244_lpi_1_dfm_1;
      operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1
          <= operator_24_14_false_AC_TRN_AC_WRAP_1_operator_24_14_false_AC_TRN_AC_WRAP_1_mux_cse_sva_1_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_4_slc_if_4_acc_1_15_svs <= 1'b0;
    end
    else if ( ~(or_dcpl_20 | or_dcpl_14 | (~((asn_sft_lpi_1_dfm_st_1[1]) & main_stage_0_2
        & if_4_for_and_mdf_sva_st_1))) ) begin
      if_4_slc_if_4_acc_1_15_svs <= if_4_acc_1_itm_15_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_4_for_and_mdf_sva_st_1 <= 1'b0;
    end
    else if ( and_dcpl_66 | or_2_tmp | (~ nand_tmp) ) begin
      if_4_for_and_mdf_sva_st_1 <= if_4_for_and_mdf_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      operator_24_14_false_AC_TRN_AC_WRAP_1_slc_operator_24_14_false_AC_TRN_AC_WRAP_1_acc_14_svs_1
          <= 1'b0;
    end
    else if ( and_dcpl_66 ) begin
      operator_24_14_false_AC_TRN_AC_WRAP_1_slc_operator_24_14_false_AC_TRN_AC_WRAP_1_acc_14_svs_1
          <= operator_24_14_false_AC_TRN_AC_WRAP_1_acc_itm_14_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      if_4_for_and_45_itm_1 <= 1'b0;
    end
    else if ( or_dcpl_1 & and_dcpl_32 & (if_4_for_mux_50_tmp[7:2]==6'b111111) & and_dcpl_25
        ) begin
      if_4_for_and_45_itm_1 <= operator_24_14_false_AC_TRN_AC_WRAP_acc_itm_14_1 &
          (~ exit_if_4_for_lpi_1_dfm_4);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      asn_sft_lpi_1_dfm_st_1 <= 10'b0000000000;
      shift_reg_1_sva_0 <= 1'b0;
    end
    else if ( or_2_tmp ) begin
      asn_sft_lpi_1_dfm_st_1 <= asn_sft_lpi_1_dfm_st_1_mx0;
      shift_reg_1_sva_0 <= shift_reg_1_sva_0_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P2_8_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1430_nl ) begin
      P2_8_1_23_10_sva <= MUX_v_14_2_2(if_4_for_1_and_52_nl, operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
          nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P2_0_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~((mux_tmp_4 | (mux_3_tmp[1]) | or_dcpl_28) & nand_tmp) ) begin
      P2_0_1_23_10_sva <= MUX_v_14_2_2(if_4_for_1_and_44_nl, operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
          nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P2_9_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1453_nl ) begin
      P2_9_1_23_10_sva <= MUX_v_14_2_2(if_4_for_1_and_53_nl, operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
          nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P2_1_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1466_nl ) begin
      P2_1_1_23_10_sva <= MUX_v_14_2_2(if_4_for_1_and_45_nl, operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
          nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P2_10_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1484_nl ) begin
      P2_10_1_23_10_sva <= MUX_v_14_2_2(if_4_for_1_and_54_nl, operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
          nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P2_2_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1510_nl ) begin
      P2_2_1_23_10_sva <= MUX_v_14_2_2(if_4_for_1_and_46_nl, operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
          nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P2_11_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1540_nl ) begin
      P2_11_1_23_10_sva <= MUX_v_14_2_2(if_4_for_1_and_55_nl, operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
          nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P2_3_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1568_nl ) begin
      P2_3_1_23_10_sva <= MUX_v_14_2_2(if_4_for_1_and_47_nl, operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
          nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P2_12_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1596_nl ) begin
      P2_12_1_23_10_sva <= MUX_v_14_2_2(if_4_for_1_and_56_nl, operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
          nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P2_4_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1625_nl ) begin
      P2_4_1_23_10_sva <= MUX_v_14_2_2(if_4_for_1_and_48_nl, operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
          nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P2_13_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1656_nl ) begin
      P2_13_1_23_10_sva <= MUX_v_14_2_2(if_4_for_1_and_57_nl, operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
          nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P2_5_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1673_nl ) begin
      P2_5_1_23_10_sva <= MUX_v_14_2_2(if_4_for_1_and_49_nl, operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
          nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P2_14_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1695_nl ) begin
      P2_14_1_23_10_sva <= MUX_v_14_2_2(if_4_for_1_and_58_nl, operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
          nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P2_6_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1718_nl ) begin
      P2_6_1_23_10_sva <= MUX_v_14_2_2(if_4_for_1_and_50_nl, operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
          nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P2_15_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( MUX_s_1_2_2(mux_1726_nl, and_258_nl, exitL_exit_approx_sva) ) begin
      P2_15_1_23_10_sva <= MUX_v_14_2_2(if_4_for_1_and_59_nl, operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
          nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P2_7_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1750_nl ) begin
      P2_7_1_23_10_sva <= MUX_v_14_2_2(if_4_for_1_and_51_nl, operator_24_14_false_AC_TRN_AC_WRAP_acc_psp_sva_1,
          nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P1_4_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1769_nl ) begin
      P1_4_1_23_10_sva <= MUX1HOT_v_14_3_2(({{13{nand_49_cse}}, nand_49_cse}), P1_4_1_23_10_sva_dfm_1_mx0,
          P1_4_1_23_10_sva_dfm_3, {nor_67_nl , nand_tmp , or_297_tmp});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P1_5_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1791_nl ) begin
      P1_5_1_23_10_sva <= MUX1HOT_v_14_3_2(({{13{nand_50_cse}}, nand_50_cse}), P1_5_1_23_10_sva_dfm_1_mx0,
          P1_5_1_23_10_sva_dfm_3, {nor_68_nl , nand_tmp , or_299_tmp});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P1_1_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1809_nl ) begin
      P1_1_1_23_10_sva <= MUX1HOT_v_14_3_2((signext_14_1(if_4_for_if_4_for_nand_4_nl)),
          P1_1_1_23_10_sva_dfm_1_mx0, P1_1_1_23_10_sva_dfm_3, {nor_69_nl , nand_tmp
          , or_301_tmp});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P1_6_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1826_nl ) begin
      P1_6_1_23_10_sva <= MUX1HOT_v_14_3_2(({{13{nand_51_cse}}, nand_51_cse}), P1_6_1_23_10_sva_dfm_1_mx0,
          P1_6_1_23_10_sva_dfm_3, {nor_70_nl , nand_tmp , or_303_tmp});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P1_2_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1845_nl ) begin
      P1_2_1_23_10_sva <= MUX1HOT_v_14_3_2((signext_14_1(if_4_for_if_4_for_nand_2_nl)),
          P1_2_1_23_10_sva_dfm_1_mx0, P1_2_1_23_10_sva_dfm_3, {nor_71_nl , nand_tmp
          , or_305_tmp});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P1_7_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( MUX_s_1_2_2(mux_1854_nl, and_263_nl, exitL_exit_approx_sva) ) begin
      P1_7_1_23_10_sva <= MUX1HOT_v_14_3_2(({{13{nand_52_cse}}, nand_52_cse}), P1_7_1_23_10_sva_dfm_1_mx0,
          P1_7_1_23_10_sva_dfm_3, {nor_72_nl , nand_tmp , or_307_tmp});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P1_3_1_23_10_sva <= 14'b00000000000000;
    end
    else if ( ~ mux_1874_nl ) begin
      P1_3_1_23_10_sva <= MUX1HOT_v_14_3_2((signext_14_1(if_4_for_if_4_for_nand_nl)),
          P1_3_1_23_10_sva_dfm_1_mx0, P1_3_1_23_10_sva_dfm_3, {nor_73_nl , nand_tmp
          , or_309_tmp});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      shift_reg_1_sva_1 <= 1'b0;
    end
    else if ( ~ nor_47_cse ) begin
      shift_reg_1_sva_1 <= shift_reg_1_sva_0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      shift_reg_1_sva_2 <= 1'b0;
    end
    else if ( ~ nor_47_cse ) begin
      shift_reg_1_sva_2 <= shift_reg_1_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      saved_reg_sva_2 <= 1'b0;
    end
    else if ( ~ or_dcpl_180 ) begin
      saved_reg_sva_2 <= shift_reg_1_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      saved_reg_sva_0 <= 1'b0;
    end
    else if ( ~ or_dcpl_180 ) begin
      saved_reg_sva_0 <= shift_reg_1_sva_0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      saved_reg_sva_1 <= 1'b0;
    end
    else if ( ~ or_dcpl_180 ) begin
      saved_reg_sva_1 <= shift_reg_1_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      reg_skip_ftd <= 1'b1;
      reg_skip_ftd_1 <= 2'b00;
    end
    else if ( skip_static_init_or_ssc ) begin
      reg_skip_ftd <= and_91_tmp_1;
      reg_skip_ftd_1 <= MUX_v_2_2_2(2'b00, skip_sva_1_1_0_1, not_402_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      or_psp <= 1'b0;
    end
    else if ( (count_sva[3:0]==4'b1111) & nand_112_cse & (count_sva[8:4]==5'b11111)
        & or_2_tmp & (count_sva[9]) ) begin
      or_psp <= or_psp_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_6 <= 1'b0;
      operator_24_14_false_AC_TRN_AC_WRAP_3_nor_m1c <= 1'b0;
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_5 <= 1'b0;
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c <= 1'b0;
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_4 <= 1'b0;
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_1 <= 1'b0;
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_3 <= 1'b0;
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_2 <= 1'b0;
    end
    else if ( operator_24_14_false_AC_TRN_AC_WRAP_3_and_38_cse ) begin
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_6 <= operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_6_mx0w0;
      operator_24_14_false_AC_TRN_AC_WRAP_3_nor_m1c <= operator_24_14_false_AC_TRN_AC_WRAP_3_nor_m1c_mx0w0;
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_5 <= operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_5_mx0w0;
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c <= operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_mx0w0;
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_4 <= operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_4_mx0w0;
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_1 <= operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_1_mx0w0;
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_3 <= operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_3_mx0w0;
      operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_2 <= operator_24_14_false_AC_TRN_AC_WRAP_3_and_m1c_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      exit_if_4_for_lpi_1_dfm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(and_298_cse, and_276_cse, or_2_tmp) ) begin
      exit_if_4_for_lpi_1_dfm <= exit_if_4_for_lpi_1_dfm_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      exit_if_4_for_lpi_1_dfm_2 <= 1'b0;
    end
    else if ( ~ nand_tmp ) begin
      exit_if_4_for_lpi_1_dfm_2 <= exit_if_4_for_lpi_1_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      j_1_3_0_lpi_1_dfm_2_2_0 <= 3'b000;
    end
    else if ( ~(mux_1306_nl | nand_tmp) ) begin
      j_1_3_0_lpi_1_dfm_2_2_0 <= j_1_3_0_sva_2[2:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      j_lpi_1_dfm_1_3_0 <= 4'b0000;
    end
    else if ( and_dcpl_67 ) begin
      j_lpi_1_dfm_1_3_0 <= if_4_for_1_acc_tmp[3:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      count_sva <= 10'b0000000000;
    end
    else if ( ~ and_dcpl_67 ) begin
      count_sva <= nl_count_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      unequal_tmp_2_1 <= 1'b0;
    end
    else if ( or_2_tmp | (~ nand_tmp) ) begin
      unequal_tmp_2_1 <= nand_tmp;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst_n ) begin
      P1_0_1_23_10_sva_rsp_0 <= 2'b00;
      P1_0_1_23_10_sva_rsp_1 <= 12'b000000000000;
    end
    else if ( mux_1772_ssc ) begin
      P1_0_1_23_10_sva_rsp_0 <= MUX_v_2_2_2(2'b00, mux_1876_nl, not_1767_nl);
      P1_0_1_23_10_sva_rsp_1 <= MUX1HOT_v_12_3_2(P1_0_1_23_10_sva_dfm_3_11_0, if_4_for_and_19_nl,
          P1_0_1_23_10_sva_dfm_1_mx0_11_0, {and_55_cse_1 , nor_cse_1 , nand_tmp});
    end
  end
  assign nl_if_4_aelse_acc_nl = conv_s2s_13_14(if_4_aelse_not_itm_1) + 14'b00000010101111;
  assign if_4_aelse_acc_nl = nl_if_4_aelse_acc_nl[13:0];
  assign if_4_for_if_4_for_or_4_nl = or_2_tmp | if_4_for_and_mdf_sva_1;
  assign or_40_nl = or_dcpl_20 | or_dcpl_14 | (~((asn_sft_lpi_1_dfm_st_1[1]) & if_4_for_and_mdf_sva_st_1));
  assign if_4_for_if_4_for_if_4_for_not_1_nl = ~ or_2_tmp;
  assign and_275_nl = (asn_sft_lpi_1_dfm_st_1==10'b1111111111) & if_4_for_and_45_itm_1;
  assign if_4_for_if_4_for_if_4_for_not_2_nl = ~ or_2_tmp;
  assign and_277_nl = (asn_sft_lpi_1_dfm_st_1==10'b1111111111) & operator_24_14_false_AC_TRN_AC_WRAP_1_slc_operator_24_14_false_AC_TRN_AC_WRAP_1_acc_14_svs_1;
  assign if_4_for_1_if_4_for_1_nand_1_nl = ~(if_4_for_1_and_stg_2_0_sva_1 & (j_lpi_1_dfm_3_0_1[3]));
  assign if_4_for_1_and_52_nl = MUX_v_14_2_2(14'b00000000000000, P2_8_1_23_10_sva_dfm_3,
      if_4_for_1_if_4_for_1_nand_1_nl);
  assign nand_91_nl = ~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_lpi_1_dfm_1_3_0==4'b1000));
  assign mux_1427_nl = MUX_s_1_2_2(mux_tmp_113, mux_tmp_96, or_325_cse);
  assign mux_1428_nl = MUX_s_1_2_2(mux_tmp_113, mux_1427_nl, or_324_cse);
  assign mux_1429_nl = MUX_s_1_2_2(nand_91_nl, mux_1428_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1419_nl = MUX_s_1_2_2(mux_tmp_105, mux_tmp_96, or_325_cse);
  assign mux_1420_nl = MUX_s_1_2_2(mux_tmp_105, mux_1419_nl, or_324_cse);
  assign mux_1430_nl = MUX_s_1_2_2(mux_1429_nl, mux_1420_nl, exitL_exit_approx_sva);
  assign if_4_for_1_if_4_for_1_nand_14_nl = ~(if_4_for_1_and_stg_2_0_sva_1 & (~ (j_lpi_1_dfm_3_0_1[3])));
  assign if_4_for_1_and_44_nl = MUX_v_14_2_2(14'b00000000000000, P2_0_1_23_10_sva_dfm_3,
      if_4_for_1_if_4_for_1_nand_14_nl);
  assign if_4_for_1_if_4_for_1_nand_3_nl = ~(if_4_for_1_and_stg_2_1_sva_1 & (j_lpi_1_dfm_3_0_1[3]));
  assign if_4_for_1_and_53_nl = MUX_v_14_2_2(14'b00000000000000, P2_9_1_23_10_sva_dfm_3,
      if_4_for_1_if_4_for_1_nand_3_nl);
  assign nand_93_nl = ~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_lpi_1_dfm_1_3_0==4'b1001));
  assign mux_1450_nl = MUX_s_1_2_2(mux_tmp_136, mux_tmp_122, or_325_cse);
  assign mux_1451_nl = MUX_s_1_2_2(mux_tmp_136, mux_1450_nl, or_324_cse);
  assign mux_1452_nl = MUX_s_1_2_2(nand_93_nl, mux_1451_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1444_nl = MUX_s_1_2_2(mux_tmp_130, mux_tmp_122, or_325_cse);
  assign mux_1445_nl = MUX_s_1_2_2(mux_tmp_130, mux_1444_nl, or_324_cse);
  assign mux_1453_nl = MUX_s_1_2_2(mux_1452_nl, mux_1445_nl, exitL_exit_approx_sva);
  assign if_4_for_1_if_4_for_1_nand_12_nl = ~(if_4_for_1_and_stg_2_1_sva_1 & (~ (j_lpi_1_dfm_3_0_1[3])));
  assign if_4_for_1_and_45_nl = MUX_v_14_2_2(14'b00000000000000, P2_1_1_23_10_sva_dfm_3,
      if_4_for_1_if_4_for_1_nand_12_nl);
  assign mux_1464_nl = MUX_s_1_2_2(or_tmp_121, mux_tmp_141, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign nand_70_nl = ~(epsilon_rsci_idat & (~ mux_tmp_141));
  assign mux_1465_nl = MUX_s_1_2_2(mux_1464_nl, nand_70_nl, exitL_exit_approx_sva);
  assign mux_1459_nl = MUX_s_1_2_2(mux_tmp_145, mux_tmp_143, or_325_cse);
  assign mux_1460_nl = MUX_s_1_2_2(mux_tmp_145, mux_1459_nl, or_324_cse);
  assign mux_1461_nl = MUX_s_1_2_2(mux_tmp_143, mux_1460_nl, first_sva);
  assign mux_1462_nl = MUX_s_1_2_2(mux_1461_nl, mux_tmp_141, epsilon_rsci_idat);
  assign mux_1463_nl = MUX_s_1_2_2(or_tmp_121, mux_1462_nl, or_2_tmp);
  assign mux_1466_nl = MUX_s_1_2_2(mux_1465_nl, mux_1463_nl, and_276_cse);
  assign if_4_for_1_if_4_for_1_nand_5_nl = ~(if_4_for_1_and_stg_2_2_sva_1 & (j_lpi_1_dfm_3_0_1[3]));
  assign if_4_for_1_and_54_nl = MUX_v_14_2_2(14'b00000000000000, P2_10_1_23_10_sva_dfm_3,
      if_4_for_1_if_4_for_1_nand_5_nl);
  assign nand_95_nl = ~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_lpi_1_dfm_1_3_0==4'b1010));
  assign mux_1481_nl = MUX_s_1_2_2(mux_tmp_167, mux_tmp_156, or_325_cse);
  assign mux_1482_nl = MUX_s_1_2_2(mux_tmp_167, mux_1481_nl, or_324_cse);
  assign mux_1483_nl = MUX_s_1_2_2(nand_95_nl, mux_1482_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1476_nl = MUX_s_1_2_2(mux_tmp_162, mux_tmp_156, or_325_cse);
  assign mux_1477_nl = MUX_s_1_2_2(mux_tmp_162, mux_1476_nl, or_324_cse);
  assign mux_1484_nl = MUX_s_1_2_2(mux_1483_nl, mux_1477_nl, exitL_exit_approx_sva);
  assign if_4_for_1_if_4_for_1_nand_10_nl = ~(if_4_for_1_and_stg_2_2_sva_1 & (~ (j_lpi_1_dfm_3_0_1[3])));
  assign if_4_for_1_and_46_nl = MUX_v_14_2_2(14'b00000000000000, P2_2_1_23_10_sva_dfm_3,
      if_4_for_1_if_4_for_1_nand_10_nl);
  assign nand_96_nl = ~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_lpi_1_dfm_1_3_0==4'b0010));
  assign mux_1500_nl = MUX_s_1_2_2(mux_tmp_186, or_tmp_143, shift_reg_1_sva_0);
  assign mux_1501_nl = MUX_s_1_2_2(mux_1500_nl, mux_tmp_173, shift_reg_1_sva_1);
  assign mux_1507_nl = MUX_s_1_2_2(mux_tmp_193, mux_1501_nl, or_325_cse);
  assign mux_1508_nl = MUX_s_1_2_2(mux_tmp_193, mux_1507_nl, or_324_cse);
  assign mux_1509_nl = MUX_s_1_2_2(nand_96_nl, mux_1508_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1488_nl = MUX_s_1_2_2(mux_tmp_174, or_tmp_143, shift_reg_1_sva_0);
  assign mux_1489_nl = MUX_s_1_2_2(mux_1488_nl, mux_tmp_173, shift_reg_1_sva_1);
  assign mux_1497_nl = MUX_s_1_2_2(mux_tmp_183, mux_1489_nl, or_325_cse);
  assign mux_1498_nl = MUX_s_1_2_2(mux_tmp_183, mux_1497_nl, or_324_cse);
  assign mux_1510_nl = MUX_s_1_2_2(mux_1509_nl, mux_1498_nl, exitL_exit_approx_sva);
  assign if_4_for_1_if_4_for_1_nand_7_nl = ~(if_4_for_1_and_stg_2_3_sva_1 & (j_lpi_1_dfm_3_0_1[3]));
  assign if_4_for_1_and_55_nl = MUX_v_14_2_2(14'b00000000000000, P2_11_1_23_10_sva_dfm_3,
      if_4_for_1_if_4_for_1_nand_7_nl);
  assign nand_98_nl = ~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_lpi_1_dfm_1_3_0==4'b1011));
  assign mux_1537_nl = MUX_s_1_2_2(not_tmp_131, mux_tmp_213, or_325_cse);
  assign mux_1538_nl = MUX_s_1_2_2(not_tmp_131, mux_1537_nl, or_324_cse);
  assign mux_1539_nl = MUX_s_1_2_2(nand_98_nl, mux_1538_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1522_nl = MUX_s_1_2_2(mux_tmp_208, mux_tmp_199, or_325_cse);
  assign mux_1523_nl = MUX_s_1_2_2(mux_tmp_208, mux_1522_nl, or_324_cse);
  assign mux_1540_nl = MUX_s_1_2_2(mux_1539_nl, mux_1523_nl, exitL_exit_approx_sva);
  assign if_4_for_1_if_4_for_1_nand_8_nl = ~(if_4_for_1_and_stg_2_3_sva_1 & (~ (j_lpi_1_dfm_3_0_1[3])));
  assign if_4_for_1_and_47_nl = MUX_v_14_2_2(14'b00000000000000, P2_3_1_23_10_sva_dfm_3,
      if_4_for_1_if_4_for_1_nand_8_nl);
  assign nand_99_nl = ~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_lpi_1_dfm_1_3_0==4'b0011));
  assign mux_1554_nl = MUX_s_1_2_2(mux_tmp_240, mux_tmp_228, shift_reg_1_sva_1);
  assign mux_1555_nl = MUX_s_1_2_2(mux_1554_nl, or_tmp_170, epsilon_rsci_idat);
  assign mux_1565_nl = MUX_s_1_2_2(mux_tmp_251, mux_1555_nl, or_325_cse);
  assign mux_1566_nl = MUX_s_1_2_2(mux_tmp_251, mux_1565_nl, or_324_cse);
  assign mux_1567_nl = MUX_s_1_2_2(nand_99_nl, mux_1566_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1542_nl = MUX_s_1_2_2(mux_tmp_228, or_tmp_170, epsilon_rsci_idat);
  assign mux_1551_nl = MUX_s_1_2_2(mux_tmp_237, mux_1542_nl, or_325_cse);
  assign mux_1552_nl = MUX_s_1_2_2(mux_tmp_237, mux_1551_nl, or_324_cse);
  assign mux_1568_nl = MUX_s_1_2_2(mux_1567_nl, mux_1552_nl, exitL_exit_approx_sva);
  assign if_4_for_1_if_4_for_1_nand_9_nl = ~(if_4_for_1_and_stg_2_4_sva_1 & (j_lpi_1_dfm_3_0_1[3]));
  assign if_4_for_1_and_56_nl = MUX_v_14_2_2(14'b00000000000000, P2_12_1_23_10_sva_dfm_3,
      if_4_for_1_if_4_for_1_nand_9_nl);
  assign or_434_nl = (~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_lpi_1_dfm_1_3_0[1:0]==2'b00)))
      | nand_101_cse;
  assign mux_1582_nl = MUX_s_1_2_2(mux_tmp_256, mux_tmp_268, shift_reg_1_sva_1);
  assign mux_1583_nl = MUX_s_1_2_2(or_tmp_190, mux_1582_nl, epsilon_rsci_idat);
  assign mux_1593_nl = MUX_s_1_2_2(mux_tmp_279, mux_1583_nl, or_325_cse);
  assign mux_1594_nl = MUX_s_1_2_2(mux_tmp_279, mux_1593_nl, or_324_cse);
  assign mux_1595_nl = MUX_s_1_2_2(or_434_nl, mux_1594_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1570_nl = MUX_s_1_2_2(or_tmp_190, mux_tmp_256, epsilon_rsci_idat);
  assign mux_1579_nl = MUX_s_1_2_2(mux_tmp_265, mux_1570_nl, or_325_cse);
  assign mux_1580_nl = MUX_s_1_2_2(mux_tmp_265, mux_1579_nl, or_324_cse);
  assign mux_1596_nl = MUX_s_1_2_2(mux_1595_nl, mux_1580_nl, exitL_exit_approx_sva);
  assign if_4_for_1_if_4_for_1_nand_6_nl = ~(if_4_for_1_and_stg_2_4_sva_1 & (~ (j_lpi_1_dfm_3_0_1[3])));
  assign if_4_for_1_and_48_nl = MUX_v_14_2_2(14'b00000000000000, P2_4_1_23_10_sva_dfm_3,
      if_4_for_1_if_4_for_1_nand_6_nl);
  assign nand_102_nl = ~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_lpi_1_dfm_1_3_0==4'b0100));
  assign mux_1622_nl = MUX_s_1_2_2(mux_tmp_308, mux_tmp_298, or_325_cse);
  assign mux_1623_nl = MUX_s_1_2_2(mux_tmp_308, mux_1622_nl, or_324_cse);
  assign mux_1624_nl = MUX_s_1_2_2(nand_102_nl, mux_1623_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1608_nl = MUX_s_1_2_2(mux_tmp_294, mux_tmp_285, or_325_cse);
  assign mux_1609_nl = MUX_s_1_2_2(mux_tmp_294, mux_1608_nl, or_324_cse);
  assign mux_1625_nl = MUX_s_1_2_2(mux_1624_nl, mux_1609_nl, exitL_exit_approx_sva);
  assign if_4_for_1_if_4_for_1_nand_11_nl = ~(if_4_for_1_and_stg_2_5_sva_1 & (j_lpi_1_dfm_3_0_1[3]));
  assign if_4_for_1_and_57_nl = MUX_v_14_2_2(14'b00000000000000, P2_13_1_23_10_sva_dfm_3,
      if_4_for_1_if_4_for_1_nand_11_nl);
  assign or_469_nl = (~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_lpi_1_dfm_1_3_0[1:0]==2'b01)))
      | nand_101_cse;
  assign mux_1644_nl = MUX_s_1_2_2(or_tmp_229, mux_tmp_330, shift_reg_1_sva_0);
  assign mux_1645_nl = MUX_s_1_2_2(mux_tmp_317, mux_1644_nl, shift_reg_1_sva_1);
  assign mux_1653_nl = MUX_s_1_2_2(mux_tmp_339, mux_1645_nl, or_325_cse);
  assign mux_1654_nl = MUX_s_1_2_2(mux_tmp_339, mux_1653_nl, or_324_cse);
  assign mux_1655_nl = MUX_s_1_2_2(or_469_nl, mux_1654_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1628_nl = MUX_s_1_2_2(or_tmp_229, mux_tmp_314, shift_reg_1_sva_0);
  assign mux_1631_nl = MUX_s_1_2_2(mux_tmp_317, mux_1628_nl, shift_reg_1_sva_1);
  assign mux_1640_nl = MUX_s_1_2_2(mux_tmp_326, mux_1631_nl, or_325_cse);
  assign mux_1641_nl = MUX_s_1_2_2(mux_tmp_326, mux_1640_nl, or_324_cse);
  assign mux_1656_nl = MUX_s_1_2_2(mux_1655_nl, mux_1641_nl, exitL_exit_approx_sva);
  assign if_4_for_1_if_4_for_1_nand_4_nl = ~(if_4_for_1_and_stg_2_5_sva_1 & (~ (j_lpi_1_dfm_3_0_1[3])));
  assign if_4_for_1_and_49_nl = MUX_v_14_2_2(14'b00000000000000, P2_5_1_23_10_sva_dfm_3,
      if_4_for_1_if_4_for_1_nand_4_nl);
  assign nand_105_nl = ~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_lpi_1_dfm_1_3_0==4'b0101));
  assign mux_1670_nl = MUX_s_1_2_2(mux_tmp_356, mux_tmp_346, or_325_cse);
  assign mux_1671_nl = MUX_s_1_2_2(mux_tmp_356, mux_1670_nl, or_324_cse);
  assign mux_1672_nl = MUX_s_1_2_2(nand_105_nl, mux_1671_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1664_nl = MUX_s_1_2_2(mux_tmp_350, mux_tmp_346, or_325_cse);
  assign mux_1665_nl = MUX_s_1_2_2(mux_tmp_350, mux_1664_nl, or_324_cse);
  assign mux_1673_nl = MUX_s_1_2_2(mux_1672_nl, mux_1665_nl, exitL_exit_approx_sva);
  assign if_4_for_1_if_4_for_1_nand_13_nl = ~(if_4_for_1_and_stg_2_6_sva_1 & (j_lpi_1_dfm_3_0_1[3]));
  assign if_4_for_1_and_58_nl = MUX_v_14_2_2(14'b00000000000000, P2_14_1_23_10_sva_dfm_3,
      if_4_for_1_if_4_for_1_nand_13_nl);
  assign or_498_nl = (~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (~ (j_lpi_1_dfm_1_3_0[0]))))
      | (j_lpi_1_dfm_1_3_0[3:1]!=3'b111);
  assign mux_1692_nl = MUX_s_1_2_2(mux_tmp_378, nand_tmp_19, or_325_cse);
  assign mux_1693_nl = MUX_s_1_2_2(mux_tmp_378, mux_1692_nl, or_324_cse);
  assign mux_1694_nl = MUX_s_1_2_2(or_498_nl, mux_1693_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1680_nl = MUX_s_1_2_2(mux_tmp_366, nand_tmp_19, or_325_cse);
  assign mux_1681_nl = MUX_s_1_2_2(mux_tmp_366, mux_1680_nl, or_324_cse);
  assign mux_1695_nl = MUX_s_1_2_2(mux_1694_nl, mux_1681_nl, exitL_exit_approx_sva);
  assign if_4_for_1_if_4_for_1_nand_2_nl = ~(if_4_for_1_and_stg_2_6_sva_1 & (~ (j_lpi_1_dfm_3_0_1[3])));
  assign if_4_for_1_and_50_nl = MUX_v_14_2_2(14'b00000000000000, P2_6_1_23_10_sva_dfm_3,
      if_4_for_1_if_4_for_1_nand_2_nl);
  assign nand_108_nl = ~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_lpi_1_dfm_1_3_0==4'b0110));
  assign mux_1715_nl = MUX_s_1_2_2(mux_tmp_401, mux_tmp_387, or_325_cse);
  assign mux_1716_nl = MUX_s_1_2_2(mux_tmp_401, mux_1715_nl, or_324_cse);
  assign mux_1717_nl = MUX_s_1_2_2(nand_108_nl, mux_1716_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1709_nl = MUX_s_1_2_2(mux_tmp_395, mux_tmp_387, or_325_cse);
  assign mux_1710_nl = MUX_s_1_2_2(mux_tmp_395, mux_1709_nl, or_324_cse);
  assign mux_1718_nl = MUX_s_1_2_2(mux_1717_nl, mux_1710_nl, exitL_exit_approx_sva);
  assign if_4_for_1_if_4_for_1_nand_15_nl = ~(if_4_for_1_and_stg_2_7_sva_1 & (j_lpi_1_dfm_3_0_1[3]));
  assign if_4_for_1_and_59_nl = MUX_v_14_2_2(14'b00000000000000, P2_15_1_23_10_sva_dfm_3,
      if_4_for_1_if_4_for_1_nand_15_nl);
  assign and_283_nl = (asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_lpi_1_dfm_1_3_0==4'b1111);
  assign and_285_nl = shift_reg_1_sva_0 & shift_reg_1_sva_1 & shift_reg_1_sva_2 &
      not_tmp_91;
  assign and_286_nl = (~((skip_sva_1_1_0_1!=2'b00) | (~ shift_reg_1_sva_0) | (~ shift_reg_1_sva_1)
      | (~ shift_reg_1_sva_2))) & not_tmp_91;
  assign mux_1724_nl = MUX_s_1_2_2(and_285_nl, and_286_nl, or_324_cse);
  assign mux_1725_nl = MUX_s_1_2_2(mux_1724_nl, mux_tmp_410, epsilon_rsci_idat);
  assign mux_1726_nl = MUX_s_1_2_2(and_283_nl, mux_1725_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign and_258_nl = epsilon_rsci_idat & mux_tmp_410;
  assign if_4_for_1_if_4_for_1_nand_nl = ~(if_4_for_1_and_stg_2_7_sva_1 & (~ (j_lpi_1_dfm_3_0_1[3])));
  assign if_4_for_1_and_51_nl = MUX_v_14_2_2(14'b00000000000000, P2_7_1_23_10_sva_dfm_3,
      if_4_for_1_if_4_for_1_nand_nl);
  assign nand_109_nl = ~((asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_lpi_1_dfm_1_3_0==4'b0111));
  assign mux_1747_nl = MUX_s_1_2_2(mux_tmp_433, mux_tmp_416, or_325_cse);
  assign mux_1748_nl = MUX_s_1_2_2(mux_tmp_433, mux_1747_nl, or_324_cse);
  assign mux_1749_nl = MUX_s_1_2_2(nand_109_nl, mux_1748_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1739_nl = MUX_s_1_2_2(mux_tmp_425, mux_tmp_416, or_325_cse);
  assign mux_1740_nl = MUX_s_1_2_2(mux_tmp_425, mux_1739_nl, or_324_cse);
  assign mux_1750_nl = MUX_s_1_2_2(mux_1749_nl, mux_1740_nl, exitL_exit_approx_sva);
  assign nor_67_nl = ~(nand_tmp | or_297_tmp);
  assign mux_1767_nl = MUX_s_1_2_2(or_tmp_310, or_546_cse, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign or_545_nl = or_dcpl_104 | or_tmp_306;
  assign mux_1768_nl = MUX_s_1_2_2(mux_1767_nl, or_545_nl, exitL_exit_approx_sva);
  assign mux_1761_nl = MUX_s_1_2_2(or_tmp_309, or_tmp_308, first_sva);
  assign mux_1759_nl = MUX_s_1_2_2(or_tmp_309, or_tmp_308, nor_149_cse);
  assign mux_1760_nl = MUX_s_1_2_2((~ mux_1759_nl), or_dcpl_100, skip_sva_1_1_0_1[1]);
  assign mux_1762_nl = MUX_s_1_2_2((~ mux_1761_nl), mux_1760_nl, or_324_cse);
  assign mux_1763_nl = MUX_s_1_2_2(mux_1762_nl, mux_tmp_440, shift_reg_1_sva_0);
  assign mux_1764_nl = MUX_s_1_2_2(mux_tmp_444, mux_1763_nl, epsilon_rsci_idat);
  assign mux_1765_nl = MUX_s_1_2_2(or_tmp_310, mux_1764_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1758_nl = MUX_s_1_2_2(mux_tmp_444, mux_tmp_440, epsilon_rsci_idat);
  assign mux_1766_nl = MUX_s_1_2_2(mux_1765_nl, mux_1758_nl, exitL_exit_approx_sva);
  assign mux_1769_nl = MUX_s_1_2_2(mux_1768_nl, mux_1766_nl, and_276_cse);
  assign nor_68_nl = ~(nand_tmp | or_299_tmp);
  assign mux_1789_nl = MUX_s_1_2_2(or_tmp_329, or_546_cse, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign or_564_nl = (~ epsilon_rsci_idat) | shift_reg_1_sva_0 | or_tmp_306;
  assign mux_1790_nl = MUX_s_1_2_2(mux_1789_nl, or_564_nl, exitL_exit_approx_sva);
  assign mux_1785_nl = MUX_s_1_2_2(or_tmp_306, (~ mux_1756_cse), shift_reg_1_sva_0);
  assign mux_1786_nl = MUX_s_1_2_2(mux_1785_nl, mux_tmp_467, epsilon_rsci_idat);
  assign mux_1787_nl = MUX_s_1_2_2(or_tmp_329, mux_1786_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign nand_110_nl = ~(shift_reg_1_sva_0 & mux_1756_cse);
  assign mux_1784_nl = MUX_s_1_2_2(nand_110_nl, mux_tmp_467, epsilon_rsci_idat);
  assign mux_1788_nl = MUX_s_1_2_2(mux_1787_nl, mux_1784_nl, exitL_exit_approx_sva);
  assign mux_1791_nl = MUX_s_1_2_2(mux_1790_nl, mux_1788_nl, and_276_cse);
  assign if_4_for_if_4_for_nand_4_nl = ~(if_4_for_and_stg_1_1_sva_1 & (~ (j_1_3_0_lpi_1_dfm_2_0_1[2])));
  assign nor_69_nl = ~(nand_tmp | or_301_tmp);
  assign nand_83_nl = ~(epsilon_rsci_idat & (~ or_tmp_334));
  assign mux_1808_nl = MUX_s_1_2_2(mux_tmp_485, nand_83_nl, exitL_exit_approx_sva);
  assign mux_1803_nl = MUX_s_1_2_2(mux_tmp_487, mux_tmp_486, first_sva);
  assign mux_1801_nl = MUX_s_1_2_2(mux_tmp_487, mux_tmp_486, nor_149_cse);
  assign mux_1802_nl = MUX_s_1_2_2(mux_1801_nl, mux_tmp_480, skip_sva_1_1_0_1[1]);
  assign mux_1804_nl = MUX_s_1_2_2(mux_1803_nl, mux_1802_nl, or_324_cse);
  assign mux_1805_nl = MUX_s_1_2_2(or_tmp_336, mux_1804_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1806_nl = MUX_s_1_2_2(mux_1805_nl, mux_tmp_485, epsilon_rsci_idat);
  assign mux_1795_nl = MUX_s_1_2_2(mux_tmp_480, mux_tmp_479, first_sva);
  assign mux_1794_nl = MUX_s_1_2_2(mux_tmp_480, mux_tmp_479, nor_159_cse);
  assign mux_1796_nl = MUX_s_1_2_2(mux_1795_nl, mux_1794_nl, or_324_cse);
  assign mux_1797_nl = MUX_s_1_2_2(mux_1796_nl, or_tmp_334, epsilon_rsci_idat);
  assign mux_1807_nl = MUX_s_1_2_2(mux_1806_nl, mux_1797_nl, exitL_exit_approx_sva);
  assign mux_1809_nl = MUX_s_1_2_2(mux_1808_nl, mux_1807_nl, and_276_cse);
  assign nor_70_nl = ~(nand_tmp | or_303_tmp);
  assign or_581_nl = epsilon_rsci_idat | or_tmp_343;
  assign mux_1825_nl = MUX_s_1_2_2(mux_tmp_509, or_581_nl, exitL_exit_approx_sva);
  assign mux_1819_nl = MUX_s_1_2_2(mux_tmp_503, or_tmp_346, first_sva);
  assign mux_1817_nl = MUX_s_1_2_2(mux_tmp_503, or_tmp_346, nor_149_cse);
  assign mux_1818_nl = MUX_s_1_2_2((~ mux_1817_nl), mux_tmp_498, skip_sva_1_1_0_1[1]);
  assign mux_1820_nl = MUX_s_1_2_2((~ mux_1819_nl), mux_1818_nl, or_324_cse);
  assign mux_1821_nl = MUX_s_1_2_2(or_tmp_347, mux_1820_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1823_nl = MUX_s_1_2_2(mux_tmp_509, mux_1821_nl, epsilon_rsci_idat);
  assign mux_1813_nl = MUX_s_1_2_2(mux_tmp_498, mux_tmp_497, first_sva);
  assign mux_1812_nl = MUX_s_1_2_2(mux_tmp_498, mux_tmp_497, nor_159_cse);
  assign mux_1814_nl = MUX_s_1_2_2(mux_1813_nl, mux_1812_nl, or_324_cse);
  assign mux_1815_nl = MUX_s_1_2_2(or_tmp_343, mux_1814_nl, epsilon_rsci_idat);
  assign mux_1824_nl = MUX_s_1_2_2(mux_1823_nl, mux_1815_nl, exitL_exit_approx_sva);
  assign mux_1826_nl = MUX_s_1_2_2(mux_1825_nl, mux_1824_nl, and_276_cse);
  assign if_4_for_if_4_for_nand_2_nl = ~(if_4_for_and_stg_1_2_sva_1 & (~ (j_1_3_0_lpi_1_dfm_2_0_1[2])));
  assign nor_71_nl = ~(nand_tmp | or_305_tmp);
  assign mux_1843_nl = MUX_s_1_2_2(or_tmp_357, nand_86_cse, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign or_608_nl = epsilon_rsci_idat | (~ shift_reg_1_sva_0) | or_tmp_356;
  assign mux_1844_nl = MUX_s_1_2_2(mux_1843_nl, or_608_nl, exitL_exit_approx_sva);
  assign mux_1839_nl = MUX_s_1_2_2(mux_1756_cse, or_tmp_356, shift_reg_1_sva_0);
  assign mux_1840_nl = MUX_s_1_2_2(mux_tmp_524, mux_1839_nl, epsilon_rsci_idat);
  assign mux_1841_nl = MUX_s_1_2_2(or_tmp_357, mux_1840_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign or_583_nl = shift_reg_1_sva_0 | mux_1756_cse;
  assign mux_1838_nl = MUX_s_1_2_2(mux_tmp_524, or_583_nl, epsilon_rsci_idat);
  assign mux_1842_nl = MUX_s_1_2_2(mux_1841_nl, mux_1838_nl, exitL_exit_approx_sva);
  assign mux_1845_nl = MUX_s_1_2_2(mux_1844_nl, mux_1842_nl, and_276_cse);
  assign nor_72_nl = ~(nand_tmp | or_307_tmp);
  assign and_293_nl = (asn_sft_lpi_1_dfm_st_1==10'b1111111111) & (j_1_3_0_lpi_1_dfm_2_2_0==3'b111)
      & (~ exit_if_4_for_lpi_1_dfm_2);
  assign mux_1853_nl = MUX_s_1_2_2(not_tmp_236, mux_tmp_538, and_294_cse);
  assign mux_1854_nl = MUX_s_1_2_2(and_293_nl, mux_1853_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1852_nl = MUX_s_1_2_2(not_tmp_236, mux_tmp_538, and_276_cse);
  assign and_263_nl = epsilon_rsci_idat & mux_1852_nl;
  assign if_4_for_if_4_for_nand_nl = ~(if_4_for_and_stg_1_3_sva_1 & (~ (j_1_3_0_lpi_1_dfm_2_0_1[2])));
  assign nor_73_nl = ~(nand_tmp | or_309_tmp);
  assign mux_1872_nl = MUX_s_1_2_2(or_tmp_370, nand_86_cse, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign nand_88_nl = ~(epsilon_rsci_idat & shift_reg_1_sva_0 & (~ or_tmp_356));
  assign mux_1873_nl = MUX_s_1_2_2(mux_1872_nl, nand_88_nl, exitL_exit_approx_sva);
  assign mux_1866_nl = MUX_s_1_2_2(nand_tmp_28, or_482_cse, first_sva);
  assign mux_1864_nl = MUX_s_1_2_2(nand_tmp_28, or_482_cse, nor_149_cse);
  assign mux_1865_nl = MUX_s_1_2_2(mux_1864_nl, nor_tmp_5, skip_sva_1_1_0_1[1]);
  assign mux_1867_nl = MUX_s_1_2_2(mux_1866_nl, mux_1865_nl, or_324_cse);
  assign mux_1868_nl = MUX_s_1_2_2(mux_tmp_549, mux_1867_nl, shift_reg_1_sva_0);
  assign mux_1869_nl = MUX_s_1_2_2((~ mux_1868_nl), mux_tmp_546, epsilon_rsci_idat);
  assign mux_1870_nl = MUX_s_1_2_2(or_tmp_370, mux_1869_nl, exitL_exit_if_4_for_2_lpi_1_dfm);
  assign mux_1863_nl = MUX_s_1_2_2((~ mux_tmp_549), mux_tmp_546, epsilon_rsci_idat);
  assign mux_1871_nl = MUX_s_1_2_2(mux_1870_nl, mux_1863_nl, exitL_exit_approx_sva);
  assign mux_1874_nl = MUX_s_1_2_2(mux_1873_nl, mux_1871_nl, and_276_cse);
  assign not_402_nl = ~ and_91_tmp_1;
  assign nor_51_nl = ~((~ exit_if_4_for_lpi_1_dfm_2) | exitL_exit_approx_sva | exitL_exit_if_4_for_2_lpi_1_dfm
      | (~ and_dcpl_66));
  assign mux_1306_nl = MUX_s_1_2_2(nor_51_nl, and_dcpl_66, j_1_3_0_sva_2[3]);
  assign nl_count_sva  = count_sva + 10'b0000000001;
  assign mux_1876_nl = MUX_v_2_2_2(P1_0_1_23_10_sva_dfm_3_13_12, P1_0_1_23_10_sva_dfm_1_mx0_13_12,
      nand_tmp);
  assign not_1767_nl = ~ nor_cse_1;
  assign if_4_for_if_4_for_nand_6_nl = ~(if_4_for_and_stg_1_0_sva_1 & (~ (j_1_3_0_lpi_1_dfm_2_0_1[2])));
  assign if_4_for_and_19_nl = MUX_v_12_2_2(12'b000000000000, P1_0_1_23_10_sva_dfm_3_11_0,
      if_4_for_if_4_for_nand_6_nl);

  function automatic [11:0] MUX1HOT_v_12_3_2;
    input [11:0] input_2;
    input [11:0] input_1;
    input [11:0] input_0;
    input [2:0] sel;
    reg [11:0] result;
  begin
    result = input_0 & {12{sel[0]}};
    result = result | (input_1 & {12{sel[1]}});
    result = result | (input_2 & {12{sel[2]}});
    MUX1HOT_v_12_3_2 = result;
  end
  endfunction


  function automatic [13:0] MUX1HOT_v_14_10_2;
    input [13:0] input_9;
    input [13:0] input_8;
    input [13:0] input_7;
    input [13:0] input_6;
    input [13:0] input_5;
    input [13:0] input_4;
    input [13:0] input_3;
    input [13:0] input_2;
    input [13:0] input_1;
    input [13:0] input_0;
    input [9:0] sel;
    reg [13:0] result;
  begin
    result = input_0 & {14{sel[0]}};
    result = result | (input_1 & {14{sel[1]}});
    result = result | (input_2 & {14{sel[2]}});
    result = result | (input_3 & {14{sel[3]}});
    result = result | (input_4 & {14{sel[4]}});
    result = result | (input_5 & {14{sel[5]}});
    result = result | (input_6 & {14{sel[6]}});
    result = result | (input_7 & {14{sel[7]}});
    result = result | (input_8 & {14{sel[8]}});
    result = result | (input_9 & {14{sel[9]}});
    MUX1HOT_v_14_10_2 = result;
  end
  endfunction


  function automatic [13:0] MUX1HOT_v_14_3_2;
    input [13:0] input_2;
    input [13:0] input_1;
    input [13:0] input_0;
    input [2:0] sel;
    reg [13:0] result;
  begin
    result = input_0 & {14{sel[0]}};
    result = result | (input_1 & {14{sel[1]}});
    result = result | (input_2 & {14{sel[2]}});
    MUX1HOT_v_14_3_2 = result;
  end
  endfunction


  function automatic [13:0] MUX1HOT_v_14_4_2;
    input [13:0] input_3;
    input [13:0] input_2;
    input [13:0] input_1;
    input [13:0] input_0;
    input [3:0] sel;
    reg [13:0] result;
  begin
    result = input_0 & {14{sel[0]}};
    result = result | (input_1 & {14{sel[1]}});
    result = result | (input_2 & {14{sel[2]}});
    result = result | (input_3 & {14{sel[3]}});
    MUX1HOT_v_14_4_2 = result;
  end
  endfunction


  function automatic [13:0] MUX1HOT_v_14_9_2;
    input [13:0] input_8;
    input [13:0] input_7;
    input [13:0] input_6;
    input [13:0] input_5;
    input [13:0] input_4;
    input [13:0] input_3;
    input [13:0] input_2;
    input [13:0] input_1;
    input [13:0] input_0;
    input [8:0] sel;
    reg [13:0] result;
  begin
    result = input_0 & {14{sel[0]}};
    result = result | (input_1 & {14{sel[1]}});
    result = result | (input_2 & {14{sel[2]}});
    result = result | (input_3 & {14{sel[3]}});
    result = result | (input_4 & {14{sel[4]}});
    result = result | (input_5 & {14{sel[5]}});
    result = result | (input_6 & {14{sel[6]}});
    result = result | (input_7 & {14{sel[7]}});
    result = result | (input_8 & {14{sel[8]}});
    MUX1HOT_v_14_9_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input  sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input  sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_16_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [13:0] input_2;
    input [13:0] input_3;
    input [13:0] input_4;
    input [13:0] input_5;
    input [13:0] input_6;
    input [13:0] input_7;
    input [13:0] input_8;
    input [13:0] input_9;
    input [13:0] input_10;
    input [13:0] input_11;
    input [13:0] input_12;
    input [13:0] input_13;
    input [13:0] input_14;
    input [13:0] input_15;
    input [3:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_14_16_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input  sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_8_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [13:0] input_2;
    input [13:0] input_3;
    input [13:0] input_4;
    input [13:0] input_5;
    input [13:0] input_6;
    input [13:0] input_7;
    input [2:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_14_8_2 = result;
  end
  endfunction


  function automatic [23:0] MUX_v_24_2_2;
    input [23:0] input_0;
    input [23:0] input_1;
    input  sel;
    reg [23:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_24_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_12_1_11;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 11;
    readslicef_12_1_11 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_13_1_12;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 12;
    readslicef_13_1_12 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_14_1_13;
    input [13:0] vector;
    reg [13:0] tmp;
  begin
    tmp = vector >> 13;
    readslicef_14_1_13 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_15_1_14;
    input [14:0] vector;
    reg [14:0] tmp;
  begin
    tmp = vector >> 14;
    readslicef_15_1_14 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_16_1_15;
    input [15:0] vector;
    reg [15:0] tmp;
  begin
    tmp = vector >> 15;
    readslicef_16_1_15 = tmp[0:0];
  end
  endfunction


  function automatic [23:0] readslicef_25_24_1;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_25_24_1 = tmp[23:0];
  end
  endfunction


  function automatic [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_7_1_6;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_7_1_6 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [13:0] signext_14_1;
    input  vector;
  begin
    signext_14_1= {{13{vector}}, vector};
  end
  endfunction


  function automatic [13:0] conv_s2s_13_14 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_14 = {vector[12], vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_15_16 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_16 = {vector[14], vector};
  end
  endfunction


  function automatic [14:0] conv_u2s_14_15 ;
    input [13:0]  vector ;
  begin
    conv_u2s_14_15 =  {1'b0, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_12 = {1'b0, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_12_13 ;
    input [11:0]  vector ;
  begin
    conv_u2u_12_13 = {1'b0, vector};
  end
  endfunction


  function automatic [13:0] conv_u2u_13_14 ;
    input [12:0]  vector ;
  begin
    conv_u2u_13_14 = {1'b0, vector};
  end
  endfunction


  function automatic [14:0] conv_u2u_14_15 ;
    input [13:0]  vector ;
  begin
    conv_u2u_14_15 = {1'b0, vector};
  end
  endfunction

endmodule



